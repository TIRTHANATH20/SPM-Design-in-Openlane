magic
tech sky130A
magscale 1 2
timestamp 1742718868
<< viali >>
rect 9965 17833 9999 17867
rect 5641 17765 5675 17799
rect 10241 17765 10275 17799
rect 4997 17629 5031 17663
rect 5365 17629 5399 17663
rect 5549 17629 5583 17663
rect 5825 17629 5859 17663
rect 8309 17629 8343 17663
rect 8769 17629 8803 17663
rect 8953 17629 8987 17663
rect 9229 17629 9263 17663
rect 9505 17629 9539 17663
rect 9689 17629 9723 17663
rect 10425 17629 10459 17663
rect 11069 17629 11103 17663
rect 12357 17629 12391 17663
rect 5089 17561 5123 17595
rect 5273 17561 5307 17595
rect 10057 17561 10091 17595
rect 5181 17493 5215 17527
rect 5457 17493 5491 17527
rect 8493 17493 8527 17527
rect 8585 17493 8619 17527
rect 9045 17493 9079 17527
rect 9413 17493 9447 17527
rect 9597 17493 9631 17527
rect 11253 17493 11287 17527
rect 12541 17493 12575 17527
rect 5917 17289 5951 17323
rect 8769 17289 8803 17323
rect 11529 17289 11563 17323
rect 1409 17153 1443 17187
rect 5457 17153 5491 17187
rect 6193 17153 6227 17187
rect 6745 17153 6779 17187
rect 9045 17153 9079 17187
rect 9597 17153 9631 17187
rect 3433 17085 3467 17119
rect 3709 17085 3743 17119
rect 5273 17085 5307 17119
rect 5549 17085 5583 17119
rect 6653 17085 6687 17119
rect 7021 17085 7055 17119
rect 7297 17085 7331 17119
rect 8861 17085 8895 17119
rect 9137 17085 9171 17119
rect 9505 17085 9539 17119
rect 9873 17085 9907 17119
rect 13001 17085 13035 17119
rect 13277 17085 13311 17119
rect 1593 16949 1627 16983
rect 5181 16949 5215 16983
rect 6009 16949 6043 16983
rect 6469 16949 6503 16983
rect 11345 16949 11379 16983
rect 5549 16745 5583 16779
rect 9229 16745 9263 16779
rect 9873 16745 9907 16779
rect 11437 16745 11471 16779
rect 6193 16609 6227 16643
rect 6469 16609 6503 16643
rect 9505 16609 9539 16643
rect 11253 16609 11287 16643
rect 1593 16541 1627 16575
rect 5089 16541 5123 16575
rect 5365 16541 5399 16575
rect 8953 16541 8987 16575
rect 9137 16541 9171 16575
rect 9229 16541 9263 16575
rect 9597 16541 9631 16575
rect 11161 16541 11195 16575
rect 1777 16405 1811 16439
rect 5181 16405 5215 16439
rect 7941 16405 7975 16439
rect 3341 16065 3375 16099
rect 3525 16065 3559 16099
rect 1409 15997 1443 16031
rect 1685 15997 1719 16031
rect 3157 15861 3191 15895
rect 3433 15861 3467 15895
rect 2789 15657 2823 15691
rect 6193 15657 6227 15691
rect 11713 15657 11747 15691
rect 1777 15589 1811 15623
rect 3893 15521 3927 15555
rect 4445 15521 4479 15555
rect 1869 15453 1903 15487
rect 2421 15453 2455 15487
rect 2973 15453 3007 15487
rect 3065 15453 3099 15487
rect 3985 15453 4019 15487
rect 7757 15453 7791 15487
rect 7849 15453 7883 15487
rect 8493 15453 8527 15487
rect 8585 15453 8619 15487
rect 9321 15453 9355 15487
rect 11621 15453 11655 15487
rect 11805 15453 11839 15487
rect 11989 15453 12023 15487
rect 12081 15453 12115 15487
rect 13093 15453 13127 15487
rect 14105 15453 14139 15487
rect 14381 15453 14415 15487
rect 14657 15453 14691 15487
rect 14749 15453 14783 15487
rect 17049 15453 17083 15487
rect 1593 15385 1627 15419
rect 2513 15385 2547 15419
rect 2697 15385 2731 15419
rect 4721 15385 4755 15419
rect 8309 15385 8343 15419
rect 9597 15385 9631 15419
rect 12265 15385 12299 15419
rect 14933 15385 14967 15419
rect 2053 15317 2087 15351
rect 2605 15317 2639 15351
rect 3433 15317 3467 15351
rect 4353 15317 4387 15351
rect 7573 15317 7607 15351
rect 8217 15317 8251 15351
rect 8585 15317 8619 15351
rect 11069 15317 11103 15351
rect 11989 15317 12023 15351
rect 13277 15317 13311 15351
rect 14197 15317 14231 15351
rect 14565 15317 14599 15351
rect 14749 15317 14783 15351
rect 16865 15317 16899 15351
rect 3525 15113 3559 15147
rect 8493 15113 8527 15147
rect 9137 15113 9171 15147
rect 15117 15113 15151 15147
rect 7021 15045 7055 15079
rect 9321 15045 9355 15079
rect 3065 14977 3099 15011
rect 3157 14977 3191 15011
rect 3341 14977 3375 15011
rect 6745 14977 6779 15011
rect 8769 14977 8803 15011
rect 9229 14977 9263 15011
rect 9413 14977 9447 15011
rect 13369 14977 13403 15011
rect 15393 14977 15427 15011
rect 8861 14909 8895 14943
rect 11529 14909 11563 14943
rect 11805 14909 11839 14943
rect 13645 14909 13679 14943
rect 15301 14909 15335 14943
rect 13277 14773 13311 14807
rect 15669 14773 15703 14807
rect 3801 14569 3835 14603
rect 7573 14569 7607 14603
rect 11897 14569 11931 14603
rect 14105 14569 14139 14603
rect 14933 14569 14967 14603
rect 17049 14569 17083 14603
rect 5549 14433 5583 14467
rect 5825 14433 5859 14467
rect 8217 14433 8251 14467
rect 10241 14433 10275 14467
rect 11621 14433 11655 14467
rect 11713 14433 11747 14467
rect 12081 14433 12115 14467
rect 14289 14433 14323 14467
rect 14749 14433 14783 14467
rect 15577 14433 15611 14467
rect 8401 14365 8435 14399
rect 8677 14365 8711 14399
rect 10149 14365 10183 14399
rect 11253 14365 11287 14399
rect 12265 14365 12299 14399
rect 12541 14365 12575 14399
rect 14381 14365 14415 14399
rect 14841 14365 14875 14399
rect 15025 14365 15059 14399
rect 15301 14365 15335 14399
rect 5273 14297 5307 14331
rect 6101 14297 6135 14331
rect 12449 14297 12483 14331
rect 8585 14229 8619 14263
rect 9781 14229 9815 14263
rect 1593 14025 1627 14059
rect 5825 14025 5859 14059
rect 10241 14025 10275 14059
rect 14749 14025 14783 14059
rect 16865 14025 16899 14059
rect 1409 13889 1443 13923
rect 5457 13889 5491 13923
rect 10241 13889 10275 13923
rect 10425 13889 10459 13923
rect 17049 13889 17083 13923
rect 5365 13821 5399 13855
rect 16497 13821 16531 13855
rect 16233 13685 16267 13719
rect 5089 13481 5123 13515
rect 1593 13413 1627 13447
rect 6745 13413 6779 13447
rect 8309 13413 8343 13447
rect 11345 13413 11379 13447
rect 5457 13345 5491 13379
rect 6101 13345 6135 13379
rect 10241 13345 10275 13379
rect 10609 13345 10643 13379
rect 1409 13277 1443 13311
rect 2881 13277 2915 13311
rect 3157 13277 3191 13311
rect 3433 13277 3467 13311
rect 3525 13277 3559 13311
rect 4997 13277 5031 13311
rect 5181 13277 5215 13311
rect 5549 13277 5583 13311
rect 5917 13277 5951 13311
rect 6285 13277 6319 13311
rect 6561 13277 6595 13311
rect 6837 13277 6871 13311
rect 6929 13277 6963 13311
rect 7665 13277 7699 13311
rect 7849 13277 7883 13311
rect 8309 13277 8343 13311
rect 8401 13277 8435 13311
rect 10149 13277 10183 13311
rect 10701 13277 10735 13311
rect 10885 13277 10919 13311
rect 11069 13277 11103 13311
rect 11161 13277 11195 13311
rect 11437 13277 11471 13311
rect 11529 13277 11563 13311
rect 12909 13277 12943 13311
rect 13185 13277 13219 13311
rect 13369 13277 13403 13311
rect 13737 13277 13771 13311
rect 17049 13277 17083 13311
rect 3249 13209 3283 13243
rect 5273 13209 5307 13243
rect 6653 13209 6687 13243
rect 8585 13209 8619 13243
rect 11253 13209 11287 13243
rect 13001 13209 13035 13243
rect 13461 13209 13495 13243
rect 13645 13209 13679 13243
rect 2697 13141 2731 13175
rect 3065 13141 3099 13175
rect 3433 13141 3467 13175
rect 6469 13141 6503 13175
rect 7665 13141 7699 13175
rect 9965 13141 9999 13175
rect 13737 13141 13771 13175
rect 16865 13141 16899 13175
rect 3157 12937 3191 12971
rect 6193 12937 6227 12971
rect 8953 12937 8987 12971
rect 11069 12937 11103 12971
rect 13277 12937 13311 12971
rect 14013 12937 14047 12971
rect 4721 12869 4755 12903
rect 9597 12869 9631 12903
rect 1409 12801 1443 12835
rect 3433 12801 3467 12835
rect 13553 12801 13587 12835
rect 14289 12801 14323 12835
rect 1685 12733 1719 12767
rect 3341 12733 3375 12767
rect 4445 12733 4479 12767
rect 7205 12733 7239 12767
rect 7481 12733 7515 12767
rect 9321 12733 9355 12767
rect 11529 12733 11563 12767
rect 11805 12733 11839 12767
rect 13369 12733 13403 12767
rect 13645 12733 13679 12767
rect 14565 12733 14599 12767
rect 3801 12665 3835 12699
rect 16037 12597 16071 12631
rect 2053 12393 2087 12427
rect 2881 12393 2915 12427
rect 5549 12393 5583 12427
rect 7481 12393 7515 12427
rect 14565 12393 14599 12427
rect 16221 12393 16255 12427
rect 8309 12325 8343 12359
rect 13369 12325 13403 12359
rect 2237 12257 2271 12291
rect 4077 12257 4111 12291
rect 7665 12257 7699 12291
rect 8125 12257 8159 12291
rect 14197 12257 14231 12291
rect 15853 12257 15887 12291
rect 16497 12257 16531 12291
rect 2329 12189 2363 12223
rect 2789 12189 2823 12223
rect 2973 12189 3007 12223
rect 3801 12189 3835 12223
rect 7757 12189 7791 12223
rect 8493 12189 8527 12223
rect 8769 12189 8803 12223
rect 13277 12189 13311 12223
rect 13461 12189 13495 12223
rect 14289 12189 14323 12223
rect 15945 12189 15979 12223
rect 16405 12189 16439 12223
rect 16589 12189 16623 12223
rect 2697 12053 2731 12087
rect 8677 12053 8711 12087
rect 10241 11849 10275 11883
rect 15117 11849 15151 11883
rect 16313 11849 16347 11883
rect 4813 11713 4847 11747
rect 4997 11713 5031 11747
rect 5733 11713 5767 11747
rect 5917 11713 5951 11747
rect 6009 11713 6043 11747
rect 7481 11713 7515 11747
rect 10057 11713 10091 11747
rect 10333 11713 10367 11747
rect 10425 11713 10459 11747
rect 10609 11713 10643 11747
rect 11529 11713 11563 11747
rect 15853 11713 15887 11747
rect 16497 11713 16531 11747
rect 16865 11713 16899 11747
rect 7573 11645 7607 11679
rect 11805 11645 11839 11679
rect 13369 11645 13403 11679
rect 13645 11645 13679 11679
rect 15761 11645 15795 11679
rect 16221 11645 16255 11679
rect 5825 11577 5859 11611
rect 4905 11509 4939 11543
rect 7205 11509 7239 11543
rect 9873 11509 9907 11543
rect 10517 11509 10551 11543
rect 13277 11509 13311 11543
rect 15577 11509 15611 11543
rect 16773 11509 16807 11543
rect 3157 11305 3191 11339
rect 6285 11305 6319 11339
rect 10701 11305 10735 11339
rect 11253 11305 11287 11339
rect 13001 11305 13035 11339
rect 3801 11237 3835 11271
rect 1409 11169 1443 11203
rect 1685 11169 1719 11203
rect 4261 11169 4295 11203
rect 4537 11169 4571 11203
rect 7205 11169 7239 11203
rect 8677 11169 8711 11203
rect 8953 11169 8987 11203
rect 10885 11169 10919 11203
rect 12817 11169 12851 11203
rect 15025 11169 15059 11203
rect 15301 11169 15335 11203
rect 16773 11169 16807 11203
rect 4169 11101 4203 11135
rect 6929 11101 6963 11135
rect 10977 11101 11011 11135
rect 12725 11101 12759 11135
rect 17049 11101 17083 11135
rect 4813 11033 4847 11067
rect 6377 11033 6411 11067
rect 6745 11033 6779 11067
rect 9229 11033 9263 11067
rect 16865 10965 16899 10999
rect 1593 10761 1627 10795
rect 2513 10761 2547 10795
rect 4353 10761 4387 10795
rect 4629 10761 4663 10795
rect 5273 10761 5307 10795
rect 7941 10761 7975 10795
rect 8217 10761 8251 10795
rect 9597 10761 9631 10795
rect 10241 10761 10275 10795
rect 10425 10761 10459 10795
rect 13001 10761 13035 10795
rect 15761 10761 15795 10795
rect 16221 10761 16255 10795
rect 2881 10693 2915 10727
rect 6009 10693 6043 10727
rect 8309 10693 8343 10727
rect 10609 10693 10643 10727
rect 16037 10693 16071 10727
rect 16497 10693 16531 10727
rect 1409 10625 1443 10659
rect 2145 10625 2179 10659
rect 2605 10625 2639 10659
rect 4905 10625 4939 10659
rect 5825 10625 5859 10659
rect 6101 10625 6135 10659
rect 7297 10625 7331 10659
rect 7757 10625 7791 10659
rect 9781 10625 9815 10659
rect 10333 10625 10367 10659
rect 10425 10625 10459 10659
rect 12357 10625 12391 10659
rect 12449 10625 12483 10659
rect 12909 10625 12943 10659
rect 13093 10625 13127 10659
rect 15577 10625 15611 10659
rect 16221 10625 16255 10659
rect 16313 10625 16347 10659
rect 17049 10625 17083 10659
rect 2237 10557 2271 10591
rect 4813 10557 4847 10591
rect 5641 10557 5675 10591
rect 9873 10557 9907 10591
rect 12817 10557 12851 10591
rect 15301 10557 15335 10591
rect 13829 10489 13863 10523
rect 16865 10489 16899 10523
rect 7573 10421 7607 10455
rect 12173 10421 12207 10455
rect 13277 10217 13311 10251
rect 15025 10217 15059 10251
rect 16129 10217 16163 10251
rect 11713 10081 11747 10115
rect 13185 10081 13219 10115
rect 15393 10081 15427 10115
rect 1409 10013 1443 10047
rect 8033 10013 8067 10047
rect 8217 10013 8251 10047
rect 11437 10013 11471 10047
rect 13461 10013 13495 10047
rect 13737 10013 13771 10047
rect 15301 10013 15335 10047
rect 16313 10013 16347 10047
rect 16589 10013 16623 10047
rect 1593 9877 1627 9911
rect 8125 9877 8159 9911
rect 13645 9877 13679 9911
rect 16497 9877 16531 9911
rect 3065 9673 3099 9707
rect 12817 9673 12851 9707
rect 15577 9673 15611 9707
rect 16405 9673 16439 9707
rect 1593 9605 1627 9639
rect 13093 9605 13127 9639
rect 1961 9537 1995 9571
rect 2697 9537 2731 9571
rect 2881 9537 2915 9571
rect 2973 9537 3007 9571
rect 3065 9537 3099 9571
rect 3249 9537 3283 9571
rect 5733 9537 5767 9571
rect 5825 9537 5859 9571
rect 6009 9537 6043 9571
rect 7849 9537 7883 9571
rect 8585 9537 8619 9571
rect 12817 9537 12851 9571
rect 12909 9537 12943 9571
rect 15577 9537 15611 9571
rect 15761 9537 15795 9571
rect 16221 9537 16255 9571
rect 16497 9537 16531 9571
rect 2053 9469 2087 9503
rect 2421 9469 2455 9503
rect 2513 9469 2547 9503
rect 7297 9469 7331 9503
rect 7573 9469 7607 9503
rect 7941 9469 7975 9503
rect 8309 9469 8343 9503
rect 8493 9469 8527 9503
rect 9137 9469 9171 9503
rect 9413 9469 9447 9503
rect 16037 9469 16071 9503
rect 8953 9401 8987 9435
rect 1501 9333 1535 9367
rect 1777 9333 1811 9367
rect 6193 9333 6227 9367
rect 7665 9333 7699 9367
rect 10885 9333 10919 9367
rect 3157 9129 3191 9163
rect 3341 9129 3375 9163
rect 8585 9129 8619 9163
rect 15853 9129 15887 9163
rect 9229 9061 9263 9095
rect 16773 9061 16807 9095
rect 1685 8993 1719 9027
rect 4077 8993 4111 9027
rect 5641 8993 5675 9027
rect 5825 8993 5859 9027
rect 6653 8993 6687 9027
rect 6929 8993 6963 9027
rect 10609 8993 10643 9027
rect 16129 8993 16163 9027
rect 16221 8993 16255 9027
rect 16589 8993 16623 9027
rect 1409 8925 1443 8959
rect 3249 8925 3283 8959
rect 3433 8925 3467 8959
rect 3525 8925 3559 8959
rect 3801 8925 3835 8959
rect 5917 8925 5951 8959
rect 6377 8925 6411 8959
rect 6561 8925 6595 8959
rect 8769 8925 8803 8959
rect 9413 8925 9447 8959
rect 10701 8925 10735 8959
rect 13093 8925 13127 8959
rect 13369 8925 13403 8959
rect 14105 8925 14139 8959
rect 16681 8925 16715 8959
rect 16865 8925 16899 8959
rect 16957 8925 16991 8959
rect 6285 8857 6319 8891
rect 8493 8857 8527 8891
rect 8677 8857 8711 8891
rect 14381 8857 14415 8891
rect 15945 8857 15979 8891
rect 5549 8789 5583 8823
rect 6469 8789 6503 8823
rect 8401 8789 8435 8823
rect 11069 8789 11103 8823
rect 1869 8585 1903 8619
rect 2973 8585 3007 8619
rect 6561 8585 6595 8619
rect 7849 8585 7883 8619
rect 10609 8585 10643 8619
rect 13921 8585 13955 8619
rect 16497 8585 16531 8619
rect 16865 8585 16899 8619
rect 4445 8517 4479 8551
rect 6377 8517 6411 8551
rect 11805 8517 11839 8551
rect 15025 8517 15059 8551
rect 1409 8449 1443 8483
rect 1685 8449 1719 8483
rect 4721 8449 4755 8483
rect 5825 8449 5859 8483
rect 6561 8449 6595 8483
rect 6653 8449 6687 8483
rect 8033 8449 8067 8483
rect 8217 8449 8251 8483
rect 8309 8449 8343 8483
rect 10057 8449 10091 8483
rect 10517 8449 10551 8483
rect 10701 8449 10735 8483
rect 13553 8449 13587 8483
rect 14749 8449 14783 8483
rect 17049 8449 17083 8483
rect 5917 8381 5951 8415
rect 9965 8381 9999 8415
rect 10425 8381 10459 8415
rect 11529 8381 11563 8415
rect 13277 8381 13311 8415
rect 13461 8381 13495 8415
rect 1593 8313 1627 8347
rect 5457 8313 5491 8347
rect 9781 8245 9815 8279
rect 1593 8041 1627 8075
rect 3341 8041 3375 8075
rect 10793 8041 10827 8075
rect 13277 8041 13311 8075
rect 9229 7905 9263 7939
rect 1409 7837 1443 7871
rect 7665 7837 7699 7871
rect 7757 7837 7791 7871
rect 8033 7837 8067 7871
rect 8217 7837 8251 7871
rect 8953 7837 8987 7871
rect 10977 7837 11011 7871
rect 11253 7837 11287 7871
rect 13185 7837 13219 7871
rect 13369 7837 13403 7871
rect 17049 7837 17083 7871
rect 3525 7769 3559 7803
rect 7941 7769 7975 7803
rect 3157 7701 3191 7735
rect 3325 7701 3359 7735
rect 7665 7701 7699 7735
rect 8217 7701 8251 7735
rect 10701 7701 10735 7735
rect 11161 7701 11195 7735
rect 16865 7701 16899 7735
rect 6193 7497 6227 7531
rect 8125 7497 8159 7531
rect 10057 7497 10091 7531
rect 13277 7497 13311 7531
rect 14013 7497 14047 7531
rect 14197 7497 14231 7531
rect 6653 7429 6687 7463
rect 10149 7429 10183 7463
rect 14105 7429 14139 7463
rect 14289 7429 14323 7463
rect 2237 7361 2271 7395
rect 2329 7361 2363 7395
rect 2513 7361 2547 7395
rect 4353 7361 4387 7395
rect 4445 7361 4479 7395
rect 8585 7361 8619 7395
rect 9873 7361 9907 7395
rect 9965 7361 9999 7395
rect 13645 7361 13679 7395
rect 14381 7361 14415 7395
rect 14565 7361 14599 7395
rect 17049 7361 17083 7395
rect 4077 7293 4111 7327
rect 4721 7293 4755 7327
rect 6377 7293 6411 7327
rect 8493 7293 8527 7327
rect 11529 7293 11563 7327
rect 11805 7293 11839 7327
rect 13369 7293 13403 7327
rect 13553 7293 13587 7327
rect 14841 7293 14875 7327
rect 2513 7225 2547 7259
rect 8217 7225 8251 7259
rect 2605 7157 2639 7191
rect 16313 7157 16347 7191
rect 16865 7157 16899 7191
rect 1672 6953 1706 6987
rect 3433 6953 3467 6987
rect 3985 6953 4019 6987
rect 7849 6953 7883 6987
rect 13369 6953 13403 6987
rect 16589 6885 16623 6919
rect 7113 6817 7147 6851
rect 7297 6817 7331 6851
rect 7757 6817 7791 6851
rect 15209 6817 15243 6851
rect 15853 6817 15887 6851
rect 1409 6749 1443 6783
rect 3249 6749 3283 6783
rect 3801 6749 3835 6783
rect 3985 6749 4019 6783
rect 5457 6749 5491 6783
rect 7389 6749 7423 6783
rect 8033 6749 8067 6783
rect 8309 6749 8343 6783
rect 13553 6749 13587 6783
rect 13829 6749 13863 6783
rect 15393 6749 15427 6783
rect 15485 6749 15519 6783
rect 16129 6749 16163 6783
rect 16405 6749 16439 6783
rect 16681 6749 16715 6783
rect 16773 6749 16807 6783
rect 4997 6681 5031 6715
rect 6193 6681 6227 6715
rect 15945 6681 15979 6715
rect 16497 6681 16531 6715
rect 3157 6613 3191 6647
rect 5089 6613 5123 6647
rect 5641 6613 5675 6647
rect 6469 6613 6503 6647
rect 8217 6613 8251 6647
rect 13737 6613 13771 6647
rect 16313 6613 16347 6647
rect 3157 6409 3191 6443
rect 11897 6409 11931 6443
rect 11161 6341 11195 6375
rect 3065 6273 3099 6307
rect 3341 6273 3375 6307
rect 8677 6273 8711 6307
rect 9229 6273 9263 6307
rect 11069 6273 11103 6307
rect 11345 6273 11379 6307
rect 11713 6273 11747 6307
rect 11989 6273 12023 6307
rect 13737 6273 13771 6307
rect 13829 6273 13863 6307
rect 14013 6273 14047 6307
rect 15761 6273 15795 6307
rect 15945 6273 15979 6307
rect 9505 6205 9539 6239
rect 10977 6205 11011 6239
rect 11069 6137 11103 6171
rect 3525 6069 3559 6103
rect 8953 6069 8987 6103
rect 11529 6069 11563 6103
rect 13921 6069 13955 6103
rect 15853 6069 15887 6103
rect 9873 5865 9907 5899
rect 13921 5865 13955 5899
rect 1593 5797 1627 5831
rect 2605 5797 2639 5831
rect 7389 5797 7423 5831
rect 9137 5797 9171 5831
rect 16865 5797 16899 5831
rect 2973 5729 3007 5763
rect 3433 5729 3467 5763
rect 3893 5729 3927 5763
rect 10057 5729 10091 5763
rect 10517 5729 10551 5763
rect 12173 5729 12207 5763
rect 15761 5729 15795 5763
rect 1409 5661 1443 5695
rect 2421 5661 2455 5695
rect 2513 5661 2547 5695
rect 3065 5661 3099 5695
rect 3985 5661 4019 5695
rect 6929 5661 6963 5695
rect 7113 5661 7147 5695
rect 7205 5661 7239 5695
rect 7573 5661 7607 5695
rect 8953 5661 8987 5695
rect 10149 5661 10183 5695
rect 10609 5661 10643 5695
rect 10793 5661 10827 5695
rect 14289 5661 14323 5695
rect 14473 5661 14507 5695
rect 14565 5661 14599 5695
rect 15669 5661 15703 5695
rect 17049 5661 17083 5695
rect 2697 5593 2731 5627
rect 7297 5593 7331 5627
rect 7481 5593 7515 5627
rect 12449 5593 12483 5627
rect 2789 5525 2823 5559
rect 4353 5525 4387 5559
rect 6745 5525 6779 5559
rect 10609 5525 10643 5559
rect 14105 5525 14139 5559
rect 16037 5525 16071 5559
rect 3525 5321 3559 5355
rect 7021 5321 7055 5355
rect 7665 5321 7699 5355
rect 9689 5321 9723 5355
rect 10885 5321 10919 5355
rect 13369 5321 13403 5355
rect 14013 5321 14047 5355
rect 16037 5321 16071 5355
rect 1869 5253 1903 5287
rect 4537 5253 4571 5287
rect 8217 5253 8251 5287
rect 11805 5253 11839 5287
rect 3433 5185 3467 5219
rect 3617 5185 3651 5219
rect 7297 5185 7331 5219
rect 10517 5185 10551 5219
rect 11529 5185 11563 5219
rect 13553 5185 13587 5219
rect 14289 5185 14323 5219
rect 1593 5117 1627 5151
rect 4261 5117 4295 5151
rect 6561 5117 6595 5151
rect 6653 5117 6687 5151
rect 7389 5117 7423 5151
rect 7941 5117 7975 5151
rect 10609 5117 10643 5151
rect 13645 5117 13679 5151
rect 14565 5117 14599 5151
rect 3341 5049 3375 5083
rect 6009 5049 6043 5083
rect 13277 5049 13311 5083
rect 6377 4981 6411 5015
rect 6837 4777 6871 4811
rect 7573 4777 7607 4811
rect 14565 4777 14599 4811
rect 5089 4641 5123 4675
rect 5365 4641 5399 4675
rect 13645 4641 13679 4675
rect 14197 4641 14231 4675
rect 16773 4641 16807 4675
rect 17049 4641 17083 4675
rect 7481 4573 7515 4607
rect 7665 4573 7699 4607
rect 13553 4573 13587 4607
rect 13737 4573 13771 4607
rect 14289 4573 14323 4607
rect 6929 4505 6963 4539
rect 7297 4505 7331 4539
rect 15301 4437 15335 4471
rect 5273 4233 5307 4267
rect 10241 4165 10275 4199
rect 5089 4097 5123 4131
rect 5365 4097 5399 4131
rect 8217 4097 8251 4131
rect 10057 4097 10091 4131
rect 12541 4097 12575 4131
rect 12725 4097 12759 4131
rect 12817 4097 12851 4131
rect 14933 4097 14967 4131
rect 15485 4097 15519 4131
rect 15577 4097 15611 4131
rect 15761 4097 15795 4131
rect 8493 4029 8527 4063
rect 15025 4029 15059 4063
rect 15669 4029 15703 4063
rect 15301 3961 15335 3995
rect 4905 3893 4939 3927
rect 9965 3893 9999 3927
rect 12357 3893 12391 3927
rect 14657 3893 14691 3927
rect 5549 3689 5583 3723
rect 7757 3689 7791 3723
rect 8953 3689 8987 3723
rect 12633 3689 12667 3723
rect 12909 3689 12943 3723
rect 16589 3689 16623 3723
rect 10333 3621 10367 3655
rect 3801 3553 3835 3587
rect 6009 3553 6043 3587
rect 9137 3553 9171 3587
rect 9689 3553 9723 3587
rect 10885 3553 10919 3587
rect 14105 3553 14139 3587
rect 15853 3553 15887 3587
rect 5917 3485 5951 3519
rect 8585 3485 8619 3519
rect 8769 3485 8803 3519
rect 9229 3485 9263 3519
rect 9597 3485 9631 3519
rect 9873 3485 9907 3519
rect 10057 3485 10091 3519
rect 10149 3485 10183 3519
rect 10425 3485 10459 3519
rect 10517 3485 10551 3519
rect 13277 3485 13311 3519
rect 13461 3485 13495 3519
rect 13553 3485 13587 3519
rect 16129 3485 16163 3519
rect 16313 3485 16347 3519
rect 16405 3485 16439 3519
rect 16773 3485 16807 3519
rect 17049 3485 17083 3519
rect 4077 3417 4111 3451
rect 5641 3417 5675 3451
rect 5825 3417 5859 3451
rect 6285 3417 6319 3451
rect 10241 3417 10275 3451
rect 11161 3417 11195 3451
rect 12817 3417 12851 3451
rect 14381 3417 14415 3451
rect 16497 3417 16531 3451
rect 16681 3417 16715 3451
rect 5917 3349 5951 3383
rect 8677 3349 8711 3383
rect 13369 3349 13403 3383
rect 15945 3349 15979 3383
rect 16865 3349 16899 3383
rect 4537 3145 4571 3179
rect 5825 3145 5859 3179
rect 8217 3145 8251 3179
rect 9045 3145 9079 3179
rect 11529 3145 11563 3179
rect 14657 3145 14691 3179
rect 15301 3145 15335 3179
rect 5181 3077 5215 3111
rect 7849 3077 7883 3111
rect 12173 3077 12207 3111
rect 14105 3077 14139 3111
rect 4721 3009 4755 3043
rect 4813 3009 4847 3043
rect 5457 3009 5491 3043
rect 5917 3009 5951 3043
rect 6101 3009 6135 3043
rect 8125 3009 8159 3043
rect 8585 3009 8619 3043
rect 10793 3009 10827 3043
rect 11713 3009 11747 3043
rect 12265 3009 12299 3043
rect 12449 3009 12483 3043
rect 14381 3009 14415 3043
rect 14841 3009 14875 3043
rect 14933 3009 14967 3043
rect 15669 3009 15703 3043
rect 17049 3009 17083 3043
rect 5365 2941 5399 2975
rect 6377 2941 6411 2975
rect 8677 2941 8711 2975
rect 10517 2941 10551 2975
rect 11805 2941 11839 2975
rect 12633 2873 12667 2907
rect 15485 2873 15519 2907
rect 16865 2873 16899 2907
rect 6009 2805 6043 2839
rect 12357 2805 12391 2839
rect 5457 2601 5491 2635
rect 7389 2601 7423 2635
rect 8493 2601 8527 2635
rect 9965 2601 9999 2635
rect 10609 2601 10643 2635
rect 11253 2601 11287 2635
rect 13185 2601 13219 2635
rect 11529 2533 11563 2567
rect 11989 2465 12023 2499
rect 5273 2397 5307 2431
rect 7205 2397 7239 2431
rect 8677 2397 8711 2431
rect 9781 2397 9815 2431
rect 10425 2397 10459 2431
rect 11069 2397 11103 2431
rect 11897 2397 11931 2431
rect 13001 2397 13035 2431
<< metal1 >>
rect 1104 17978 17388 18000
rect 1104 17926 2985 17978
rect 3037 17926 3049 17978
rect 3101 17926 3113 17978
rect 3165 17926 3177 17978
rect 3229 17926 3241 17978
rect 3293 17926 7056 17978
rect 7108 17926 7120 17978
rect 7172 17926 7184 17978
rect 7236 17926 7248 17978
rect 7300 17926 7312 17978
rect 7364 17926 11127 17978
rect 11179 17926 11191 17978
rect 11243 17926 11255 17978
rect 11307 17926 11319 17978
rect 11371 17926 11383 17978
rect 11435 17926 15198 17978
rect 15250 17926 15262 17978
rect 15314 17926 15326 17978
rect 15378 17926 15390 17978
rect 15442 17926 15454 17978
rect 15506 17926 17388 17978
rect 1104 17904 17388 17926
rect 9582 17824 9588 17876
rect 9640 17864 9646 17876
rect 9953 17867 10011 17873
rect 9953 17864 9965 17867
rect 9640 17836 9965 17864
rect 9640 17824 9646 17836
rect 9953 17833 9965 17836
rect 9999 17864 10011 17867
rect 12342 17864 12348 17876
rect 9999 17836 12348 17864
rect 9999 17833 10011 17836
rect 9953 17827 10011 17833
rect 12342 17824 12348 17836
rect 12400 17824 12406 17876
rect 5074 17756 5080 17808
rect 5132 17796 5138 17808
rect 5629 17799 5687 17805
rect 5629 17796 5641 17799
rect 5132 17768 5641 17796
rect 5132 17756 5138 17768
rect 5629 17765 5641 17768
rect 5675 17765 5687 17799
rect 5629 17759 5687 17765
rect 8938 17756 8944 17808
rect 8996 17796 9002 17808
rect 10229 17799 10287 17805
rect 10229 17796 10241 17799
rect 8996 17768 10241 17796
rect 8996 17756 9002 17768
rect 10229 17765 10241 17768
rect 10275 17765 10287 17799
rect 10229 17759 10287 17765
rect 5166 17688 5172 17740
rect 5224 17728 5230 17740
rect 9030 17728 9036 17740
rect 5224 17700 5856 17728
rect 5224 17688 5230 17700
rect 4062 17620 4068 17672
rect 4120 17660 4126 17672
rect 4985 17663 5043 17669
rect 4985 17660 4997 17663
rect 4120 17632 4997 17660
rect 4120 17620 4126 17632
rect 4985 17629 4997 17632
rect 5031 17629 5043 17663
rect 4985 17623 5043 17629
rect 5353 17663 5411 17669
rect 5353 17629 5365 17663
rect 5399 17660 5411 17663
rect 5442 17660 5448 17672
rect 5399 17632 5448 17660
rect 5399 17629 5411 17632
rect 5353 17623 5411 17629
rect 5442 17620 5448 17632
rect 5500 17620 5506 17672
rect 5828 17669 5856 17700
rect 8772 17700 9036 17728
rect 5537 17663 5595 17669
rect 5537 17629 5549 17663
rect 5583 17629 5595 17663
rect 5537 17623 5595 17629
rect 5813 17663 5871 17669
rect 5813 17629 5825 17663
rect 5859 17629 5871 17663
rect 5813 17623 5871 17629
rect 8297 17663 8355 17669
rect 8297 17629 8309 17663
rect 8343 17660 8355 17663
rect 8386 17660 8392 17672
rect 8343 17632 8392 17660
rect 8343 17629 8355 17632
rect 8297 17623 8355 17629
rect 5074 17552 5080 17604
rect 5132 17552 5138 17604
rect 5258 17552 5264 17604
rect 5316 17552 5322 17604
rect 5552 17592 5580 17623
rect 8386 17620 8392 17632
rect 8444 17620 8450 17672
rect 8772 17669 8800 17700
rect 9030 17688 9036 17700
rect 9088 17688 9094 17740
rect 9398 17688 9404 17740
rect 9456 17728 9462 17740
rect 9456 17700 9720 17728
rect 9456 17688 9462 17700
rect 8757 17663 8815 17669
rect 8757 17629 8769 17663
rect 8803 17629 8815 17663
rect 8757 17623 8815 17629
rect 8938 17620 8944 17672
rect 8996 17620 9002 17672
rect 9122 17620 9128 17672
rect 9180 17660 9186 17672
rect 9692 17669 9720 17700
rect 9217 17663 9275 17669
rect 9217 17660 9229 17663
rect 9180 17632 9229 17660
rect 9180 17620 9186 17632
rect 9217 17629 9229 17632
rect 9263 17629 9275 17663
rect 9217 17623 9275 17629
rect 9493 17663 9551 17669
rect 9493 17629 9505 17663
rect 9539 17629 9551 17663
rect 9493 17623 9551 17629
rect 9677 17663 9735 17669
rect 9677 17629 9689 17663
rect 9723 17629 9735 17663
rect 9677 17623 9735 17629
rect 5902 17592 5908 17604
rect 5368 17564 5908 17592
rect 5169 17527 5227 17533
rect 5169 17493 5181 17527
rect 5215 17524 5227 17527
rect 5368 17524 5396 17564
rect 5902 17552 5908 17564
rect 5960 17552 5966 17604
rect 9508 17592 9536 17623
rect 9766 17620 9772 17672
rect 9824 17660 9830 17672
rect 10413 17663 10471 17669
rect 10413 17660 10425 17663
rect 9824 17632 10425 17660
rect 9824 17620 9830 17632
rect 10413 17629 10425 17632
rect 10459 17629 10471 17663
rect 10413 17623 10471 17629
rect 10962 17620 10968 17672
rect 11020 17660 11026 17672
rect 11057 17663 11115 17669
rect 11057 17660 11069 17663
rect 11020 17632 11069 17660
rect 11020 17620 11026 17632
rect 11057 17629 11069 17632
rect 11103 17629 11115 17663
rect 11057 17623 11115 17629
rect 12250 17620 12256 17672
rect 12308 17660 12314 17672
rect 12345 17663 12403 17669
rect 12345 17660 12357 17663
rect 12308 17632 12357 17660
rect 12308 17620 12314 17632
rect 12345 17629 12357 17632
rect 12391 17629 12403 17663
rect 12345 17623 12403 17629
rect 9232 17564 9536 17592
rect 9232 17536 9260 17564
rect 10042 17552 10048 17604
rect 10100 17592 10106 17604
rect 13078 17592 13084 17604
rect 10100 17564 13084 17592
rect 10100 17552 10106 17564
rect 13078 17552 13084 17564
rect 13136 17552 13142 17604
rect 5215 17496 5396 17524
rect 5445 17527 5503 17533
rect 5215 17493 5227 17496
rect 5169 17487 5227 17493
rect 5445 17493 5457 17527
rect 5491 17524 5503 17527
rect 5534 17524 5540 17536
rect 5491 17496 5540 17524
rect 5491 17493 5503 17496
rect 5445 17487 5503 17493
rect 5534 17484 5540 17496
rect 5592 17484 5598 17536
rect 8478 17484 8484 17536
rect 8536 17484 8542 17536
rect 8570 17484 8576 17536
rect 8628 17484 8634 17536
rect 8662 17484 8668 17536
rect 8720 17524 8726 17536
rect 9033 17527 9091 17533
rect 9033 17524 9045 17527
rect 8720 17496 9045 17524
rect 8720 17484 8726 17496
rect 9033 17493 9045 17496
rect 9079 17493 9091 17527
rect 9033 17487 9091 17493
rect 9214 17484 9220 17536
rect 9272 17484 9278 17536
rect 9398 17484 9404 17536
rect 9456 17484 9462 17536
rect 9490 17484 9496 17536
rect 9548 17524 9554 17536
rect 9585 17527 9643 17533
rect 9585 17524 9597 17527
rect 9548 17496 9597 17524
rect 9548 17484 9554 17496
rect 9585 17493 9597 17496
rect 9631 17493 9643 17527
rect 9585 17487 9643 17493
rect 11241 17527 11299 17533
rect 11241 17493 11253 17527
rect 11287 17524 11299 17527
rect 11514 17524 11520 17536
rect 11287 17496 11520 17524
rect 11287 17493 11299 17496
rect 11241 17487 11299 17493
rect 11514 17484 11520 17496
rect 11572 17484 11578 17536
rect 12526 17484 12532 17536
rect 12584 17484 12590 17536
rect 1104 17434 17388 17456
rect 1104 17382 3645 17434
rect 3697 17382 3709 17434
rect 3761 17382 3773 17434
rect 3825 17382 3837 17434
rect 3889 17382 3901 17434
rect 3953 17382 7716 17434
rect 7768 17382 7780 17434
rect 7832 17382 7844 17434
rect 7896 17382 7908 17434
rect 7960 17382 7972 17434
rect 8024 17382 11787 17434
rect 11839 17382 11851 17434
rect 11903 17382 11915 17434
rect 11967 17382 11979 17434
rect 12031 17382 12043 17434
rect 12095 17382 15858 17434
rect 15910 17382 15922 17434
rect 15974 17382 15986 17434
rect 16038 17382 16050 17434
rect 16102 17382 16114 17434
rect 16166 17382 17388 17434
rect 1104 17360 17388 17382
rect 5902 17280 5908 17332
rect 5960 17280 5966 17332
rect 8757 17323 8815 17329
rect 8757 17289 8769 17323
rect 8803 17320 8815 17323
rect 8938 17320 8944 17332
rect 8803 17292 8944 17320
rect 8803 17289 8815 17292
rect 8757 17283 8815 17289
rect 8938 17280 8944 17292
rect 8996 17320 9002 17332
rect 9122 17320 9128 17332
rect 8996 17292 9128 17320
rect 8996 17280 9002 17292
rect 9122 17280 9128 17292
rect 9180 17280 9186 17332
rect 9306 17320 9312 17332
rect 9232 17292 9312 17320
rect 4154 17212 4160 17264
rect 4212 17212 4218 17264
rect 5534 17212 5540 17264
rect 5592 17252 5598 17264
rect 9232 17252 9260 17292
rect 9306 17280 9312 17292
rect 9364 17320 9370 17332
rect 11517 17323 11575 17329
rect 11517 17320 11529 17323
rect 9364 17292 11529 17320
rect 9364 17280 9370 17292
rect 11517 17289 11529 17292
rect 11563 17289 11575 17323
rect 11517 17283 11575 17289
rect 5592 17224 6684 17252
rect 5592 17212 5598 17224
rect 842 17144 848 17196
rect 900 17184 906 17196
rect 1397 17187 1455 17193
rect 1397 17184 1409 17187
rect 900 17156 1409 17184
rect 900 17144 906 17156
rect 1397 17153 1409 17156
rect 1443 17153 1455 17187
rect 1397 17147 1455 17153
rect 5442 17144 5448 17196
rect 5500 17144 5506 17196
rect 5994 17144 6000 17196
rect 6052 17184 6058 17196
rect 6181 17187 6239 17193
rect 6181 17184 6193 17187
rect 6052 17156 6193 17184
rect 6052 17144 6058 17156
rect 6181 17153 6193 17156
rect 6227 17153 6239 17187
rect 6181 17147 6239 17153
rect 3418 17076 3424 17128
rect 3476 17076 3482 17128
rect 3697 17119 3755 17125
rect 3697 17085 3709 17119
rect 3743 17116 3755 17119
rect 5261 17119 5319 17125
rect 5261 17116 5273 17119
rect 3743 17088 5273 17116
rect 3743 17085 3755 17088
rect 3697 17079 3755 17085
rect 5261 17085 5273 17088
rect 5307 17085 5319 17119
rect 5261 17079 5319 17085
rect 5537 17119 5595 17125
rect 5537 17085 5549 17119
rect 5583 17116 5595 17119
rect 6270 17116 6276 17128
rect 5583 17088 6276 17116
rect 5583 17085 5595 17088
rect 5537 17079 5595 17085
rect 6270 17076 6276 17088
rect 6328 17116 6334 17128
rect 6546 17116 6552 17128
rect 6328 17088 6552 17116
rect 6328 17076 6334 17088
rect 6546 17076 6552 17088
rect 6604 17076 6610 17128
rect 6656 17125 6684 17224
rect 8956 17224 9260 17252
rect 6730 17144 6736 17196
rect 6788 17144 6794 17196
rect 8386 17144 8392 17196
rect 8444 17144 8450 17196
rect 6641 17119 6699 17125
rect 6641 17085 6653 17119
rect 6687 17085 6699 17119
rect 7009 17119 7067 17125
rect 7009 17116 7021 17119
rect 6641 17079 6699 17085
rect 6886 17088 7021 17116
rect 6886 17048 6914 17088
rect 7009 17085 7021 17088
rect 7055 17085 7067 17119
rect 7009 17079 7067 17085
rect 7285 17119 7343 17125
rect 7285 17085 7297 17119
rect 7331 17116 7343 17119
rect 8849 17119 8907 17125
rect 8849 17116 8861 17119
rect 7331 17088 8861 17116
rect 7331 17085 7343 17088
rect 7285 17079 7343 17085
rect 8849 17085 8861 17088
rect 8895 17085 8907 17119
rect 8956 17116 8984 17224
rect 9033 17187 9091 17193
rect 9033 17153 9045 17187
rect 9079 17184 9091 17187
rect 9398 17184 9404 17196
rect 9079 17156 9404 17184
rect 9079 17153 9091 17156
rect 9033 17147 9091 17153
rect 9398 17144 9404 17156
rect 9456 17144 9462 17196
rect 9582 17144 9588 17196
rect 9640 17144 9646 17196
rect 9125 17119 9183 17125
rect 9125 17116 9137 17119
rect 8956 17088 9137 17116
rect 8849 17079 8907 17085
rect 9125 17085 9137 17088
rect 9171 17085 9183 17119
rect 9125 17079 9183 17085
rect 9214 17076 9220 17128
rect 9272 17116 9278 17128
rect 9493 17119 9551 17125
rect 9493 17116 9505 17119
rect 9272 17088 9505 17116
rect 9272 17076 9278 17088
rect 9493 17085 9505 17088
rect 9539 17085 9551 17119
rect 9493 17079 9551 17085
rect 9858 17076 9864 17128
rect 9916 17076 9922 17128
rect 10870 17076 10876 17128
rect 10928 17116 10934 17128
rect 10980 17116 11008 17170
rect 11900 17116 11928 17170
rect 10928 17088 11928 17116
rect 10928 17076 10934 17088
rect 12986 17076 12992 17128
rect 13044 17076 13050 17128
rect 13265 17119 13323 17125
rect 13265 17085 13277 17119
rect 13311 17085 13323 17119
rect 13265 17079 13323 17085
rect 6104 17020 6914 17048
rect 6104 16992 6132 17020
rect 1578 16940 1584 16992
rect 1636 16940 1642 16992
rect 5169 16983 5227 16989
rect 5169 16949 5181 16983
rect 5215 16980 5227 16983
rect 5258 16980 5264 16992
rect 5215 16952 5264 16980
rect 5215 16949 5227 16952
rect 5169 16943 5227 16949
rect 5258 16940 5264 16952
rect 5316 16940 5322 16992
rect 5997 16983 6055 16989
rect 5997 16949 6009 16983
rect 6043 16980 6055 16983
rect 6086 16980 6092 16992
rect 6043 16952 6092 16980
rect 6043 16949 6055 16952
rect 5997 16943 6055 16949
rect 6086 16940 6092 16952
rect 6144 16940 6150 16992
rect 6454 16940 6460 16992
rect 6512 16940 6518 16992
rect 9122 16940 9128 16992
rect 9180 16980 9186 16992
rect 9582 16980 9588 16992
rect 9180 16952 9588 16980
rect 9180 16940 9186 16952
rect 9582 16940 9588 16952
rect 9640 16940 9646 16992
rect 10318 16940 10324 16992
rect 10376 16980 10382 16992
rect 11333 16983 11391 16989
rect 11333 16980 11345 16983
rect 10376 16952 11345 16980
rect 10376 16940 10382 16952
rect 11333 16949 11345 16952
rect 11379 16949 11391 16983
rect 11333 16943 11391 16949
rect 12342 16940 12348 16992
rect 12400 16980 12406 16992
rect 13280 16980 13308 17079
rect 12400 16952 13308 16980
rect 12400 16940 12406 16952
rect 1104 16890 17388 16912
rect 1104 16838 2985 16890
rect 3037 16838 3049 16890
rect 3101 16838 3113 16890
rect 3165 16838 3177 16890
rect 3229 16838 3241 16890
rect 3293 16838 7056 16890
rect 7108 16838 7120 16890
rect 7172 16838 7184 16890
rect 7236 16838 7248 16890
rect 7300 16838 7312 16890
rect 7364 16838 11127 16890
rect 11179 16838 11191 16890
rect 11243 16838 11255 16890
rect 11307 16838 11319 16890
rect 11371 16838 11383 16890
rect 11435 16838 15198 16890
rect 15250 16838 15262 16890
rect 15314 16838 15326 16890
rect 15378 16838 15390 16890
rect 15442 16838 15454 16890
rect 15506 16838 17388 16890
rect 1104 16816 17388 16838
rect 5442 16736 5448 16788
rect 5500 16776 5506 16788
rect 5537 16779 5595 16785
rect 5537 16776 5549 16779
rect 5500 16748 5549 16776
rect 5500 16736 5506 16748
rect 5537 16745 5549 16748
rect 5583 16745 5595 16779
rect 5537 16739 5595 16745
rect 5994 16736 6000 16788
rect 6052 16776 6058 16788
rect 6052 16748 9168 16776
rect 6052 16736 6058 16748
rect 9140 16708 9168 16748
rect 9214 16736 9220 16788
rect 9272 16736 9278 16788
rect 9858 16736 9864 16788
rect 9916 16736 9922 16788
rect 11425 16779 11483 16785
rect 11425 16745 11437 16779
rect 11471 16776 11483 16779
rect 12986 16776 12992 16788
rect 11471 16748 12992 16776
rect 11471 16745 11483 16748
rect 11425 16739 11483 16745
rect 12986 16736 12992 16748
rect 13044 16736 13050 16788
rect 10042 16708 10048 16720
rect 9140 16680 10048 16708
rect 10042 16668 10048 16680
rect 10100 16668 10106 16720
rect 6086 16600 6092 16652
rect 6144 16640 6150 16652
rect 6181 16643 6239 16649
rect 6181 16640 6193 16643
rect 6144 16612 6193 16640
rect 6144 16600 6150 16612
rect 6181 16609 6193 16612
rect 6227 16609 6239 16643
rect 6181 16603 6239 16609
rect 6454 16600 6460 16652
rect 6512 16600 6518 16652
rect 9490 16600 9496 16652
rect 9548 16600 9554 16652
rect 11241 16643 11299 16649
rect 11241 16609 11253 16643
rect 11287 16640 11299 16643
rect 11698 16640 11704 16652
rect 11287 16612 11704 16640
rect 11287 16609 11299 16612
rect 11241 16603 11299 16609
rect 11698 16600 11704 16612
rect 11756 16600 11762 16652
rect 1578 16532 1584 16584
rect 1636 16532 1642 16584
rect 5074 16532 5080 16584
rect 5132 16532 5138 16584
rect 5258 16532 5264 16584
rect 5316 16572 5322 16584
rect 5353 16575 5411 16581
rect 5353 16572 5365 16575
rect 5316 16544 5365 16572
rect 5316 16532 5322 16544
rect 5353 16541 5365 16544
rect 5399 16541 5411 16575
rect 8386 16572 8392 16584
rect 7590 16544 8392 16572
rect 5353 16535 5411 16541
rect 8386 16532 8392 16544
rect 8444 16532 8450 16584
rect 8938 16532 8944 16584
rect 8996 16532 9002 16584
rect 9030 16532 9036 16584
rect 9088 16572 9094 16584
rect 9125 16575 9183 16581
rect 9125 16572 9137 16575
rect 9088 16544 9137 16572
rect 9088 16532 9094 16544
rect 9125 16541 9137 16544
rect 9171 16541 9183 16575
rect 9125 16535 9183 16541
rect 9217 16575 9275 16581
rect 9217 16541 9229 16575
rect 9263 16541 9275 16575
rect 9217 16535 9275 16541
rect 5994 16504 6000 16516
rect 1780 16476 6000 16504
rect 1578 16396 1584 16448
rect 1636 16436 1642 16448
rect 1780 16445 1808 16476
rect 5994 16464 6000 16476
rect 6052 16464 6058 16516
rect 8202 16464 8208 16516
rect 8260 16504 8266 16516
rect 9232 16504 9260 16535
rect 9306 16532 9312 16584
rect 9364 16572 9370 16584
rect 9585 16575 9643 16581
rect 9585 16572 9597 16575
rect 9364 16544 9597 16572
rect 9364 16532 9370 16544
rect 9585 16541 9597 16544
rect 9631 16541 9643 16575
rect 9585 16535 9643 16541
rect 11149 16575 11207 16581
rect 11149 16541 11161 16575
rect 11195 16572 11207 16575
rect 11606 16572 11612 16584
rect 11195 16544 11612 16572
rect 11195 16541 11207 16544
rect 11149 16535 11207 16541
rect 11606 16532 11612 16544
rect 11664 16532 11670 16584
rect 8260 16476 9260 16504
rect 8260 16464 8266 16476
rect 1765 16439 1823 16445
rect 1765 16436 1777 16439
rect 1636 16408 1777 16436
rect 1636 16396 1642 16408
rect 1765 16405 1777 16408
rect 1811 16405 1823 16439
rect 1765 16399 1823 16405
rect 5074 16396 5080 16448
rect 5132 16436 5138 16448
rect 5169 16439 5227 16445
rect 5169 16436 5181 16439
rect 5132 16408 5181 16436
rect 5132 16396 5138 16408
rect 5169 16405 5181 16408
rect 5215 16405 5227 16439
rect 5169 16399 5227 16405
rect 7929 16439 7987 16445
rect 7929 16405 7941 16439
rect 7975 16436 7987 16439
rect 8110 16436 8116 16448
rect 7975 16408 8116 16436
rect 7975 16405 7987 16408
rect 7929 16399 7987 16405
rect 8110 16396 8116 16408
rect 8168 16396 8174 16448
rect 1104 16346 17388 16368
rect 1104 16294 3645 16346
rect 3697 16294 3709 16346
rect 3761 16294 3773 16346
rect 3825 16294 3837 16346
rect 3889 16294 3901 16346
rect 3953 16294 7716 16346
rect 7768 16294 7780 16346
rect 7832 16294 7844 16346
rect 7896 16294 7908 16346
rect 7960 16294 7972 16346
rect 8024 16294 11787 16346
rect 11839 16294 11851 16346
rect 11903 16294 11915 16346
rect 11967 16294 11979 16346
rect 12031 16294 12043 16346
rect 12095 16294 15858 16346
rect 15910 16294 15922 16346
rect 15974 16294 15986 16346
rect 16038 16294 16050 16346
rect 16102 16294 16114 16346
rect 16166 16294 17388 16346
rect 1104 16272 17388 16294
rect 4154 16164 4160 16176
rect 2898 16136 4160 16164
rect 4154 16124 4160 16136
rect 4212 16164 4218 16176
rect 5166 16164 5172 16176
rect 4212 16136 5172 16164
rect 4212 16124 4218 16136
rect 5166 16124 5172 16136
rect 5224 16124 5230 16176
rect 3326 16056 3332 16108
rect 3384 16056 3390 16108
rect 3510 16056 3516 16108
rect 3568 16056 3574 16108
rect 1394 15988 1400 16040
rect 1452 15988 1458 16040
rect 1670 15988 1676 16040
rect 1728 15988 1734 16040
rect 2774 15852 2780 15904
rect 2832 15892 2838 15904
rect 3145 15895 3203 15901
rect 3145 15892 3157 15895
rect 2832 15864 3157 15892
rect 2832 15852 2838 15864
rect 3145 15861 3157 15864
rect 3191 15861 3203 15895
rect 3145 15855 3203 15861
rect 3421 15895 3479 15901
rect 3421 15861 3433 15895
rect 3467 15892 3479 15895
rect 3878 15892 3884 15904
rect 3467 15864 3884 15892
rect 3467 15861 3479 15864
rect 3421 15855 3479 15861
rect 3878 15852 3884 15864
rect 3936 15852 3942 15904
rect 1104 15802 17388 15824
rect 1104 15750 2985 15802
rect 3037 15750 3049 15802
rect 3101 15750 3113 15802
rect 3165 15750 3177 15802
rect 3229 15750 3241 15802
rect 3293 15750 7056 15802
rect 7108 15750 7120 15802
rect 7172 15750 7184 15802
rect 7236 15750 7248 15802
rect 7300 15750 7312 15802
rect 7364 15750 11127 15802
rect 11179 15750 11191 15802
rect 11243 15750 11255 15802
rect 11307 15750 11319 15802
rect 11371 15750 11383 15802
rect 11435 15750 15198 15802
rect 15250 15750 15262 15802
rect 15314 15750 15326 15802
rect 15378 15750 15390 15802
rect 15442 15750 15454 15802
rect 15506 15750 17388 15802
rect 1104 15728 17388 15750
rect 1670 15648 1676 15700
rect 1728 15688 1734 15700
rect 2777 15691 2835 15697
rect 2777 15688 2789 15691
rect 1728 15660 2789 15688
rect 1728 15648 1734 15660
rect 2777 15657 2789 15660
rect 2823 15657 2835 15691
rect 2777 15651 2835 15657
rect 3234 15648 3240 15700
rect 3292 15688 3298 15700
rect 4062 15688 4068 15700
rect 3292 15660 4068 15688
rect 3292 15648 3298 15660
rect 4062 15648 4068 15660
rect 4120 15688 4126 15700
rect 6181 15691 6239 15697
rect 4120 15660 6132 15688
rect 4120 15648 4126 15660
rect 1394 15580 1400 15632
rect 1452 15620 1458 15632
rect 1765 15623 1823 15629
rect 1765 15620 1777 15623
rect 1452 15592 1777 15620
rect 1452 15580 1458 15592
rect 1765 15589 1777 15592
rect 1811 15620 1823 15623
rect 3418 15620 3424 15632
rect 1811 15592 3424 15620
rect 1811 15589 1823 15592
rect 1765 15583 1823 15589
rect 3418 15580 3424 15592
rect 3476 15620 3482 15632
rect 6104 15620 6132 15660
rect 6181 15657 6193 15691
rect 6227 15688 6239 15691
rect 6270 15688 6276 15700
rect 6227 15660 6276 15688
rect 6227 15657 6239 15660
rect 6181 15651 6239 15657
rect 6270 15648 6276 15660
rect 6328 15648 6334 15700
rect 11698 15648 11704 15700
rect 11756 15648 11762 15700
rect 12618 15620 12624 15632
rect 3476 15592 4476 15620
rect 6104 15592 6914 15620
rect 3476 15580 3482 15592
rect 3234 15552 3240 15564
rect 2424 15524 3240 15552
rect 1026 15444 1032 15496
rect 1084 15484 1090 15496
rect 2424 15493 2452 15524
rect 3234 15512 3240 15524
rect 3292 15512 3298 15564
rect 3878 15512 3884 15564
rect 3936 15512 3942 15564
rect 4448 15561 4476 15592
rect 4433 15555 4491 15561
rect 4433 15521 4445 15555
rect 4479 15552 4491 15555
rect 5258 15552 5264 15564
rect 4479 15524 5264 15552
rect 4479 15521 4491 15524
rect 4433 15515 4491 15521
rect 5258 15512 5264 15524
rect 5316 15512 5322 15564
rect 6886 15552 6914 15592
rect 11992 15592 12624 15620
rect 8202 15552 8208 15564
rect 6886 15524 8208 15552
rect 8202 15512 8208 15524
rect 8260 15552 8266 15564
rect 8260 15524 8616 15552
rect 8260 15512 8266 15524
rect 1857 15487 1915 15493
rect 1857 15484 1869 15487
rect 1084 15456 1869 15484
rect 1084 15444 1090 15456
rect 1857 15453 1869 15456
rect 1903 15453 1915 15487
rect 1857 15447 1915 15453
rect 2409 15487 2467 15493
rect 2409 15453 2421 15487
rect 2455 15453 2467 15487
rect 2866 15484 2872 15496
rect 2409 15447 2467 15453
rect 2516 15456 2872 15484
rect 1578 15376 1584 15428
rect 1636 15376 1642 15428
rect 2516 15425 2544 15456
rect 2866 15444 2872 15456
rect 2924 15444 2930 15496
rect 2958 15444 2964 15496
rect 3016 15444 3022 15496
rect 3053 15487 3111 15493
rect 3053 15453 3065 15487
rect 3099 15484 3111 15487
rect 3970 15484 3976 15496
rect 3099 15456 3976 15484
rect 3099 15453 3111 15456
rect 3053 15447 3111 15453
rect 3970 15444 3976 15456
rect 4028 15444 4034 15496
rect 7558 15444 7564 15496
rect 7616 15484 7622 15496
rect 7745 15487 7803 15493
rect 7745 15484 7757 15487
rect 7616 15456 7757 15484
rect 7616 15444 7622 15456
rect 7745 15453 7757 15456
rect 7791 15453 7803 15487
rect 7745 15447 7803 15453
rect 7837 15487 7895 15493
rect 7837 15453 7849 15487
rect 7883 15453 7895 15487
rect 7837 15447 7895 15453
rect 2501 15419 2559 15425
rect 2501 15416 2513 15419
rect 2056 15388 2513 15416
rect 2056 15357 2084 15388
rect 2501 15385 2513 15388
rect 2547 15385 2559 15419
rect 2501 15379 2559 15385
rect 2682 15376 2688 15428
rect 2740 15376 2746 15428
rect 4709 15419 4767 15425
rect 4709 15385 4721 15419
rect 4755 15385 4767 15419
rect 4709 15379 4767 15385
rect 2041 15351 2099 15357
rect 2041 15317 2053 15351
rect 2087 15317 2099 15351
rect 2041 15311 2099 15317
rect 2593 15351 2651 15357
rect 2593 15317 2605 15351
rect 2639 15348 2651 15351
rect 3326 15348 3332 15360
rect 2639 15320 3332 15348
rect 2639 15317 2651 15320
rect 2593 15311 2651 15317
rect 3326 15308 3332 15320
rect 3384 15348 3390 15360
rect 3421 15351 3479 15357
rect 3421 15348 3433 15351
rect 3384 15320 3433 15348
rect 3384 15308 3390 15320
rect 3421 15317 3433 15320
rect 3467 15317 3479 15351
rect 3421 15311 3479 15317
rect 4341 15351 4399 15357
rect 4341 15317 4353 15351
rect 4387 15348 4399 15351
rect 4724 15348 4752 15379
rect 5166 15376 5172 15428
rect 5224 15376 5230 15428
rect 7466 15376 7472 15428
rect 7524 15416 7530 15428
rect 7852 15416 7880 15447
rect 8478 15444 8484 15496
rect 8536 15444 8542 15496
rect 8588 15493 8616 15524
rect 8573 15487 8631 15493
rect 8573 15453 8585 15487
rect 8619 15453 8631 15487
rect 8573 15447 8631 15453
rect 9306 15444 9312 15496
rect 9364 15444 9370 15496
rect 11609 15487 11667 15493
rect 11609 15453 11621 15487
rect 11655 15453 11667 15487
rect 11609 15447 11667 15453
rect 7524 15388 7880 15416
rect 7524 15376 7530 15388
rect 8294 15376 8300 15428
rect 8352 15376 8358 15428
rect 9582 15376 9588 15428
rect 9640 15376 9646 15428
rect 10870 15416 10876 15428
rect 10810 15388 10876 15416
rect 10870 15376 10876 15388
rect 10928 15376 10934 15428
rect 11624 15416 11652 15447
rect 11698 15444 11704 15496
rect 11756 15484 11762 15496
rect 11992 15493 12020 15592
rect 12618 15580 12624 15592
rect 12676 15620 12682 15632
rect 12676 15592 13308 15620
rect 12676 15580 12682 15592
rect 11793 15487 11851 15493
rect 11793 15484 11805 15487
rect 11756 15456 11805 15484
rect 11756 15444 11762 15456
rect 11793 15453 11805 15456
rect 11839 15453 11851 15487
rect 11793 15447 11851 15453
rect 11977 15487 12035 15493
rect 11977 15453 11989 15487
rect 12023 15453 12035 15487
rect 11977 15447 12035 15453
rect 12069 15487 12127 15493
rect 12069 15453 12081 15487
rect 12115 15484 12127 15487
rect 12526 15484 12532 15496
rect 12115 15456 12532 15484
rect 12115 15453 12127 15456
rect 12069 15447 12127 15453
rect 12526 15444 12532 15456
rect 12584 15444 12590 15496
rect 13078 15444 13084 15496
rect 13136 15444 13142 15496
rect 11624 15388 12020 15416
rect 4387 15320 4752 15348
rect 4387 15317 4399 15320
rect 4341 15311 4399 15317
rect 7006 15308 7012 15360
rect 7064 15348 7070 15360
rect 7561 15351 7619 15357
rect 7561 15348 7573 15351
rect 7064 15320 7573 15348
rect 7064 15308 7070 15320
rect 7561 15317 7573 15320
rect 7607 15317 7619 15351
rect 7561 15311 7619 15317
rect 8205 15351 8263 15357
rect 8205 15317 8217 15351
rect 8251 15348 8263 15351
rect 8573 15351 8631 15357
rect 8573 15348 8585 15351
rect 8251 15320 8585 15348
rect 8251 15317 8263 15320
rect 8205 15311 8263 15317
rect 8573 15317 8585 15320
rect 8619 15348 8631 15351
rect 9398 15348 9404 15360
rect 8619 15320 9404 15348
rect 8619 15317 8631 15320
rect 8573 15311 8631 15317
rect 9398 15308 9404 15320
rect 9456 15308 9462 15360
rect 11057 15351 11115 15357
rect 11057 15317 11069 15351
rect 11103 15348 11115 15351
rect 11606 15348 11612 15360
rect 11103 15320 11612 15348
rect 11103 15317 11115 15320
rect 11057 15311 11115 15317
rect 11606 15308 11612 15320
rect 11664 15308 11670 15360
rect 11992 15357 12020 15388
rect 12250 15376 12256 15428
rect 12308 15376 12314 15428
rect 13280 15416 13308 15592
rect 14108 15592 15056 15620
rect 14108 15493 14136 15592
rect 14918 15552 14924 15564
rect 14384 15524 14924 15552
rect 14384 15493 14412 15524
rect 14918 15512 14924 15524
rect 14976 15512 14982 15564
rect 14093 15487 14151 15493
rect 14093 15453 14105 15487
rect 14139 15453 14151 15487
rect 14093 15447 14151 15453
rect 14369 15487 14427 15493
rect 14369 15453 14381 15487
rect 14415 15453 14427 15487
rect 14369 15447 14427 15453
rect 14645 15487 14703 15493
rect 14645 15453 14657 15487
rect 14691 15453 14703 15487
rect 14645 15447 14703 15453
rect 14737 15487 14795 15493
rect 14737 15453 14749 15487
rect 14783 15484 14795 15487
rect 15028 15484 15056 15592
rect 16574 15484 16580 15496
rect 14783 15456 16580 15484
rect 14783 15453 14795 15456
rect 14737 15447 14795 15453
rect 14660 15416 14688 15447
rect 16574 15444 16580 15456
rect 16632 15444 16638 15496
rect 17034 15444 17040 15496
rect 17092 15444 17098 15496
rect 13280 15388 14688 15416
rect 14918 15376 14924 15428
rect 14976 15376 14982 15428
rect 11977 15351 12035 15357
rect 11977 15317 11989 15351
rect 12023 15348 12035 15351
rect 12158 15348 12164 15360
rect 12023 15320 12164 15348
rect 12023 15317 12035 15320
rect 11977 15311 12035 15317
rect 12158 15308 12164 15320
rect 12216 15308 12222 15360
rect 13262 15308 13268 15360
rect 13320 15308 13326 15360
rect 14182 15308 14188 15360
rect 14240 15308 14246 15360
rect 14550 15308 14556 15360
rect 14608 15308 14614 15360
rect 14734 15308 14740 15360
rect 14792 15308 14798 15360
rect 16850 15308 16856 15360
rect 16908 15308 16914 15360
rect 1104 15258 17388 15280
rect 1104 15206 3645 15258
rect 3697 15206 3709 15258
rect 3761 15206 3773 15258
rect 3825 15206 3837 15258
rect 3889 15206 3901 15258
rect 3953 15206 7716 15258
rect 7768 15206 7780 15258
rect 7832 15206 7844 15258
rect 7896 15206 7908 15258
rect 7960 15206 7972 15258
rect 8024 15206 11787 15258
rect 11839 15206 11851 15258
rect 11903 15206 11915 15258
rect 11967 15206 11979 15258
rect 12031 15206 12043 15258
rect 12095 15206 15858 15258
rect 15910 15206 15922 15258
rect 15974 15206 15986 15258
rect 16038 15206 16050 15258
rect 16102 15206 16114 15258
rect 16166 15206 17388 15258
rect 1104 15184 17388 15206
rect 2958 15104 2964 15156
rect 3016 15144 3022 15156
rect 3510 15144 3516 15156
rect 3016 15116 3516 15144
rect 3016 15104 3022 15116
rect 3510 15104 3516 15116
rect 3568 15104 3574 15156
rect 8294 15104 8300 15156
rect 8352 15144 8358 15156
rect 8481 15147 8539 15153
rect 8481 15144 8493 15147
rect 8352 15116 8493 15144
rect 8352 15104 8358 15116
rect 8481 15113 8493 15116
rect 8527 15113 8539 15147
rect 8481 15107 8539 15113
rect 9125 15147 9183 15153
rect 9125 15113 9137 15147
rect 9171 15144 9183 15147
rect 9582 15144 9588 15156
rect 9171 15116 9588 15144
rect 9171 15113 9183 15116
rect 9125 15107 9183 15113
rect 9582 15104 9588 15116
rect 9640 15104 9646 15156
rect 14918 15104 14924 15156
rect 14976 15144 14982 15156
rect 15105 15147 15163 15153
rect 15105 15144 15117 15147
rect 14976 15116 15117 15144
rect 14976 15104 14982 15116
rect 15105 15113 15117 15116
rect 15151 15113 15163 15147
rect 15105 15107 15163 15113
rect 2774 15036 2780 15088
rect 2832 15076 2838 15088
rect 2832 15048 3372 15076
rect 2832 15036 2838 15048
rect 2866 14968 2872 15020
rect 2924 15008 2930 15020
rect 3344 15017 3372 15048
rect 7006 15036 7012 15088
rect 7064 15036 7070 15088
rect 8386 15076 8392 15088
rect 8234 15048 8392 15076
rect 8386 15036 8392 15048
rect 8444 15036 8450 15088
rect 9309 15079 9367 15085
rect 9309 15076 9321 15079
rect 8864 15048 9321 15076
rect 3053 15011 3111 15017
rect 3053 15008 3065 15011
rect 2924 14980 3065 15008
rect 2924 14968 2930 14980
rect 3053 14977 3065 14980
rect 3099 14977 3111 15011
rect 3053 14971 3111 14977
rect 3145 15011 3203 15017
rect 3145 14977 3157 15011
rect 3191 14977 3203 15011
rect 3145 14971 3203 14977
rect 3329 15011 3387 15017
rect 3329 14977 3341 15011
rect 3375 14977 3387 15011
rect 3329 14971 3387 14977
rect 3160 14940 3188 14971
rect 6086 14968 6092 15020
rect 6144 15008 6150 15020
rect 6733 15011 6791 15017
rect 6733 15008 6745 15011
rect 6144 14980 6745 15008
rect 6144 14968 6150 14980
rect 6733 14977 6745 14980
rect 6779 14977 6791 15011
rect 6733 14971 6791 14977
rect 8757 15011 8815 15017
rect 8757 14977 8769 15011
rect 8803 14977 8815 15011
rect 8757 14971 8815 14977
rect 3510 14940 3516 14952
rect 3160 14912 3516 14940
rect 3510 14900 3516 14912
rect 3568 14940 3574 14952
rect 5074 14940 5080 14952
rect 3568 14912 5080 14940
rect 3568 14900 3574 14912
rect 5074 14900 5080 14912
rect 5132 14900 5138 14952
rect 7466 14900 7472 14952
rect 7524 14940 7530 14952
rect 8772 14940 8800 14971
rect 8864 14949 8892 15048
rect 9309 15045 9321 15048
rect 9355 15045 9367 15079
rect 15654 15076 15660 15088
rect 14858 15048 15660 15076
rect 9309 15039 9367 15045
rect 15654 15036 15660 15048
rect 15712 15036 15718 15088
rect 9217 15011 9275 15017
rect 9217 15008 9229 15011
rect 8956 14980 9229 15008
rect 7524 14912 8800 14940
rect 8849 14943 8907 14949
rect 7524 14900 7530 14912
rect 8849 14909 8861 14943
rect 8895 14909 8907 14943
rect 8849 14903 8907 14909
rect 5092 14804 5120 14900
rect 7374 14804 7380 14816
rect 5092 14776 7380 14804
rect 7374 14764 7380 14776
rect 7432 14764 7438 14816
rect 7558 14764 7564 14816
rect 7616 14804 7622 14816
rect 8956 14804 8984 14980
rect 9217 14977 9229 14980
rect 9263 14977 9275 15011
rect 9217 14971 9275 14977
rect 9398 14968 9404 15020
rect 9456 14968 9462 15020
rect 12894 14968 12900 15020
rect 12952 14968 12958 15020
rect 13262 14968 13268 15020
rect 13320 15008 13326 15020
rect 13357 15011 13415 15017
rect 13357 15008 13369 15011
rect 13320 14980 13369 15008
rect 13320 14968 13326 14980
rect 13357 14977 13369 14980
rect 13403 14977 13415 15011
rect 15381 15011 15439 15017
rect 15381 15008 15393 15011
rect 13357 14971 13415 14977
rect 14844 14980 15393 15008
rect 11517 14943 11575 14949
rect 11517 14909 11529 14943
rect 11563 14909 11575 14943
rect 11517 14903 11575 14909
rect 11793 14943 11851 14949
rect 11793 14909 11805 14943
rect 11839 14940 11851 14943
rect 11882 14940 11888 14952
rect 11839 14912 11888 14940
rect 11839 14909 11851 14912
rect 11793 14903 11851 14909
rect 7616 14776 8984 14804
rect 11532 14804 11560 14903
rect 11882 14900 11888 14912
rect 11940 14900 11946 14952
rect 13633 14943 13691 14949
rect 13633 14909 13645 14943
rect 13679 14940 13691 14943
rect 14090 14940 14096 14952
rect 13679 14912 14096 14940
rect 13679 14909 13691 14912
rect 13633 14903 13691 14909
rect 14090 14900 14096 14912
rect 14148 14900 14154 14952
rect 14366 14900 14372 14952
rect 14424 14940 14430 14952
rect 14844 14940 14872 14980
rect 15381 14977 15393 14980
rect 15427 14977 15439 15011
rect 15381 14971 15439 14977
rect 14424 14912 14872 14940
rect 14424 14900 14430 14912
rect 14918 14900 14924 14952
rect 14976 14940 14982 14952
rect 15289 14943 15347 14949
rect 15289 14940 15301 14943
rect 14976 14912 15301 14940
rect 14976 14900 14982 14912
rect 15289 14909 15301 14912
rect 15335 14909 15347 14943
rect 15289 14903 15347 14909
rect 11790 14804 11796 14816
rect 11532 14776 11796 14804
rect 7616 14764 7622 14776
rect 11790 14764 11796 14776
rect 11848 14764 11854 14816
rect 12250 14764 12256 14816
rect 12308 14804 12314 14816
rect 13265 14807 13323 14813
rect 13265 14804 13277 14807
rect 12308 14776 13277 14804
rect 12308 14764 12314 14776
rect 13265 14773 13277 14776
rect 13311 14773 13323 14807
rect 13265 14767 13323 14773
rect 15562 14764 15568 14816
rect 15620 14804 15626 14816
rect 15657 14807 15715 14813
rect 15657 14804 15669 14807
rect 15620 14776 15669 14804
rect 15620 14764 15626 14776
rect 15657 14773 15669 14776
rect 15703 14773 15715 14807
rect 15657 14767 15715 14773
rect 1104 14714 17388 14736
rect 1104 14662 2985 14714
rect 3037 14662 3049 14714
rect 3101 14662 3113 14714
rect 3165 14662 3177 14714
rect 3229 14662 3241 14714
rect 3293 14662 7056 14714
rect 7108 14662 7120 14714
rect 7172 14662 7184 14714
rect 7236 14662 7248 14714
rect 7300 14662 7312 14714
rect 7364 14662 11127 14714
rect 11179 14662 11191 14714
rect 11243 14662 11255 14714
rect 11307 14662 11319 14714
rect 11371 14662 11383 14714
rect 11435 14662 15198 14714
rect 15250 14662 15262 14714
rect 15314 14662 15326 14714
rect 15378 14662 15390 14714
rect 15442 14662 15454 14714
rect 15506 14662 17388 14714
rect 1104 14640 17388 14662
rect 3789 14603 3847 14609
rect 3789 14569 3801 14603
rect 3835 14600 3847 14603
rect 3970 14600 3976 14612
rect 3835 14572 3976 14600
rect 3835 14569 3847 14572
rect 3789 14563 3847 14569
rect 3970 14560 3976 14572
rect 4028 14560 4034 14612
rect 7466 14560 7472 14612
rect 7524 14600 7530 14612
rect 7561 14603 7619 14609
rect 7561 14600 7573 14603
rect 7524 14572 7573 14600
rect 7524 14560 7530 14572
rect 7561 14569 7573 14572
rect 7607 14569 7619 14603
rect 7561 14563 7619 14569
rect 11882 14560 11888 14612
rect 11940 14560 11946 14612
rect 14090 14560 14096 14612
rect 14148 14560 14154 14612
rect 14918 14560 14924 14612
rect 14976 14560 14982 14612
rect 17034 14560 17040 14612
rect 17092 14560 17098 14612
rect 7374 14492 7380 14544
rect 7432 14532 7438 14544
rect 8662 14532 8668 14544
rect 7432 14504 8668 14532
rect 7432 14492 7438 14504
rect 8662 14492 8668 14504
rect 8720 14492 8726 14544
rect 11790 14492 11796 14544
rect 11848 14532 11854 14544
rect 12342 14532 12348 14544
rect 11848 14504 12348 14532
rect 11848 14492 11854 14504
rect 12342 14492 12348 14504
rect 12400 14492 12406 14544
rect 14568 14504 15056 14532
rect 14568 14476 14596 14504
rect 5258 14424 5264 14476
rect 5316 14464 5322 14476
rect 5537 14467 5595 14473
rect 5537 14464 5549 14467
rect 5316 14436 5549 14464
rect 5316 14424 5322 14436
rect 5537 14433 5549 14436
rect 5583 14433 5595 14467
rect 5537 14427 5595 14433
rect 5813 14467 5871 14473
rect 5813 14433 5825 14467
rect 5859 14464 5871 14467
rect 6086 14464 6092 14476
rect 5859 14436 6092 14464
rect 5859 14433 5871 14436
rect 5813 14427 5871 14433
rect 6086 14424 6092 14436
rect 6144 14424 6150 14476
rect 7558 14424 7564 14476
rect 7616 14464 7622 14476
rect 8205 14467 8263 14473
rect 8205 14464 8217 14467
rect 7616 14436 8217 14464
rect 7616 14424 7622 14436
rect 8205 14433 8217 14436
rect 8251 14433 8263 14467
rect 8205 14427 8263 14433
rect 10226 14424 10232 14476
rect 10284 14424 10290 14476
rect 11606 14424 11612 14476
rect 11664 14424 11670 14476
rect 11698 14424 11704 14476
rect 11756 14464 11762 14476
rect 12069 14467 12127 14473
rect 12069 14464 12081 14467
rect 11756 14436 12081 14464
rect 11756 14424 11762 14436
rect 12069 14433 12081 14436
rect 12115 14433 12127 14467
rect 12069 14427 12127 14433
rect 14277 14467 14335 14473
rect 14277 14433 14289 14467
rect 14323 14464 14335 14467
rect 14550 14464 14556 14476
rect 14323 14436 14556 14464
rect 14323 14433 14335 14436
rect 14277 14427 14335 14433
rect 14550 14424 14556 14436
rect 14608 14424 14614 14476
rect 14734 14424 14740 14476
rect 14792 14424 14798 14476
rect 7668 14368 7972 14396
rect 5166 14328 5172 14340
rect 4830 14300 5172 14328
rect 5166 14288 5172 14300
rect 5224 14288 5230 14340
rect 5261 14331 5319 14337
rect 5261 14297 5273 14331
rect 5307 14297 5319 14331
rect 5261 14291 5319 14297
rect 5276 14260 5304 14291
rect 6086 14288 6092 14340
rect 6144 14288 6150 14340
rect 7558 14328 7564 14340
rect 7314 14300 7564 14328
rect 7558 14288 7564 14300
rect 7616 14288 7622 14340
rect 7668 14260 7696 14368
rect 7944 14328 7972 14368
rect 8294 14356 8300 14408
rect 8352 14396 8358 14408
rect 8389 14399 8447 14405
rect 8389 14396 8401 14399
rect 8352 14368 8401 14396
rect 8352 14356 8358 14368
rect 8389 14365 8401 14368
rect 8435 14365 8447 14399
rect 8389 14359 8447 14365
rect 8478 14356 8484 14408
rect 8536 14396 8542 14408
rect 8665 14399 8723 14405
rect 8665 14396 8677 14399
rect 8536 14368 8677 14396
rect 8536 14356 8542 14368
rect 8665 14365 8677 14368
rect 8711 14365 8723 14399
rect 8665 14359 8723 14365
rect 10137 14399 10195 14405
rect 10137 14365 10149 14399
rect 10183 14396 10195 14399
rect 10318 14396 10324 14408
rect 10183 14368 10324 14396
rect 10183 14365 10195 14368
rect 10137 14359 10195 14365
rect 10318 14356 10324 14368
rect 10376 14356 10382 14408
rect 11241 14399 11299 14405
rect 11241 14365 11253 14399
rect 11287 14396 11299 14399
rect 12158 14396 12164 14408
rect 11287 14368 12164 14396
rect 11287 14365 11299 14368
rect 11241 14359 11299 14365
rect 12158 14356 12164 14368
rect 12216 14356 12222 14408
rect 12250 14356 12256 14408
rect 12308 14356 12314 14408
rect 12526 14356 12532 14408
rect 12584 14356 12590 14408
rect 13262 14356 13268 14408
rect 13320 14396 13326 14408
rect 13320 14368 14320 14396
rect 13320 14356 13326 14368
rect 14292 14340 14320 14368
rect 14366 14356 14372 14408
rect 14424 14356 14430 14408
rect 14752 14396 14780 14424
rect 15028 14405 15056 14504
rect 15562 14424 15568 14476
rect 15620 14424 15626 14476
rect 14829 14399 14887 14405
rect 14829 14396 14841 14399
rect 14752 14368 14841 14396
rect 14829 14365 14841 14368
rect 14875 14365 14887 14399
rect 14829 14359 14887 14365
rect 15013 14399 15071 14405
rect 15013 14365 15025 14399
rect 15059 14365 15071 14399
rect 15013 14359 15071 14365
rect 15289 14399 15347 14405
rect 15289 14365 15301 14399
rect 15335 14365 15347 14399
rect 15289 14359 15347 14365
rect 7944 14300 9812 14328
rect 5276 14232 7696 14260
rect 8573 14263 8631 14269
rect 8573 14229 8585 14263
rect 8619 14260 8631 14263
rect 8662 14260 8668 14272
rect 8619 14232 8668 14260
rect 8619 14229 8631 14232
rect 8573 14223 8631 14229
rect 8662 14220 8668 14232
rect 8720 14220 8726 14272
rect 9784 14269 9812 14300
rect 12434 14288 12440 14340
rect 12492 14328 12498 14340
rect 14182 14328 14188 14340
rect 12492 14300 14188 14328
rect 12492 14288 12498 14300
rect 14182 14288 14188 14300
rect 14240 14288 14246 14340
rect 14274 14288 14280 14340
rect 14332 14328 14338 14340
rect 15304 14328 15332 14359
rect 14332 14300 15332 14328
rect 14332 14288 14338 14300
rect 15654 14288 15660 14340
rect 15712 14328 15718 14340
rect 15712 14300 16054 14328
rect 15712 14288 15718 14300
rect 9769 14263 9827 14269
rect 9769 14229 9781 14263
rect 9815 14229 9827 14263
rect 9769 14223 9827 14229
rect 1104 14170 17388 14192
rect 1104 14118 3645 14170
rect 3697 14118 3709 14170
rect 3761 14118 3773 14170
rect 3825 14118 3837 14170
rect 3889 14118 3901 14170
rect 3953 14118 7716 14170
rect 7768 14118 7780 14170
rect 7832 14118 7844 14170
rect 7896 14118 7908 14170
rect 7960 14118 7972 14170
rect 8024 14118 11787 14170
rect 11839 14118 11851 14170
rect 11903 14118 11915 14170
rect 11967 14118 11979 14170
rect 12031 14118 12043 14170
rect 12095 14118 15858 14170
rect 15910 14118 15922 14170
rect 15974 14118 15986 14170
rect 16038 14118 16050 14170
rect 16102 14118 16114 14170
rect 16166 14118 17388 14170
rect 1104 14096 17388 14118
rect 1581 14059 1639 14065
rect 1581 14025 1593 14059
rect 1627 14056 1639 14059
rect 2774 14056 2780 14068
rect 1627 14028 2780 14056
rect 1627 14025 1639 14028
rect 1581 14019 1639 14025
rect 2774 14016 2780 14028
rect 2832 14016 2838 14068
rect 5813 14059 5871 14065
rect 5813 14025 5825 14059
rect 5859 14056 5871 14059
rect 6086 14056 6092 14068
rect 5859 14028 6092 14056
rect 5859 14025 5871 14028
rect 5813 14019 5871 14025
rect 6086 14016 6092 14028
rect 6144 14016 6150 14068
rect 7558 14016 7564 14068
rect 7616 14056 7622 14068
rect 8386 14056 8392 14068
rect 7616 14028 8392 14056
rect 7616 14016 7622 14028
rect 8386 14016 8392 14028
rect 8444 14016 8450 14068
rect 10226 14016 10232 14068
rect 10284 14016 10290 14068
rect 14366 14016 14372 14068
rect 14424 14056 14430 14068
rect 14737 14059 14795 14065
rect 14737 14056 14749 14059
rect 14424 14028 14749 14056
rect 14424 14016 14430 14028
rect 14737 14025 14749 14028
rect 14783 14025 14795 14059
rect 14737 14019 14795 14025
rect 16574 14016 16580 14068
rect 16632 14056 16638 14068
rect 16853 14059 16911 14065
rect 16853 14056 16865 14059
rect 16632 14028 16865 14056
rect 16632 14016 16638 14028
rect 16853 14025 16865 14028
rect 16899 14025 16911 14059
rect 16853 14019 16911 14025
rect 15654 13948 15660 14000
rect 15712 13948 15718 14000
rect 1394 13880 1400 13932
rect 1452 13880 1458 13932
rect 5445 13923 5503 13929
rect 5445 13889 5457 13923
rect 5491 13920 5503 13923
rect 5534 13920 5540 13932
rect 5491 13892 5540 13920
rect 5491 13889 5503 13892
rect 5445 13883 5503 13889
rect 5534 13880 5540 13892
rect 5592 13880 5598 13932
rect 10134 13880 10140 13932
rect 10192 13920 10198 13932
rect 10229 13923 10287 13929
rect 10229 13920 10241 13923
rect 10192 13892 10241 13920
rect 10192 13880 10198 13892
rect 10229 13889 10241 13892
rect 10275 13889 10287 13923
rect 10229 13883 10287 13889
rect 10410 13880 10416 13932
rect 10468 13880 10474 13932
rect 17034 13880 17040 13932
rect 17092 13880 17098 13932
rect 5350 13812 5356 13864
rect 5408 13812 5414 13864
rect 14274 13812 14280 13864
rect 14332 13852 14338 13864
rect 16485 13855 16543 13861
rect 16485 13852 16497 13855
rect 14332 13824 16497 13852
rect 14332 13812 14338 13824
rect 16485 13821 16497 13824
rect 16531 13821 16543 13855
rect 16485 13815 16543 13821
rect 16206 13676 16212 13728
rect 16264 13725 16270 13728
rect 16264 13719 16279 13725
rect 16267 13685 16279 13719
rect 16264 13679 16279 13685
rect 16264 13676 16270 13679
rect 1104 13626 17388 13648
rect 1104 13574 2985 13626
rect 3037 13574 3049 13626
rect 3101 13574 3113 13626
rect 3165 13574 3177 13626
rect 3229 13574 3241 13626
rect 3293 13574 7056 13626
rect 7108 13574 7120 13626
rect 7172 13574 7184 13626
rect 7236 13574 7248 13626
rect 7300 13574 7312 13626
rect 7364 13574 11127 13626
rect 11179 13574 11191 13626
rect 11243 13574 11255 13626
rect 11307 13574 11319 13626
rect 11371 13574 11383 13626
rect 11435 13574 15198 13626
rect 15250 13574 15262 13626
rect 15314 13574 15326 13626
rect 15378 13574 15390 13626
rect 15442 13574 15454 13626
rect 15506 13574 17388 13626
rect 1104 13552 17388 13574
rect 5077 13515 5135 13521
rect 5077 13481 5089 13515
rect 5123 13512 5135 13515
rect 5350 13512 5356 13524
rect 5123 13484 5356 13512
rect 5123 13481 5135 13484
rect 5077 13475 5135 13481
rect 5350 13472 5356 13484
rect 5408 13472 5414 13524
rect 1581 13447 1639 13453
rect 1581 13413 1593 13447
rect 1627 13444 1639 13447
rect 6733 13447 6791 13453
rect 6733 13444 6745 13447
rect 1627 13416 4660 13444
rect 1627 13413 1639 13416
rect 1581 13407 1639 13413
rect 2774 13336 2780 13388
rect 2832 13376 2838 13388
rect 2832 13348 3188 13376
rect 2832 13336 2838 13348
rect 842 13268 848 13320
rect 900 13308 906 13320
rect 3160 13317 3188 13348
rect 3326 13336 3332 13388
rect 3384 13376 3390 13388
rect 3384 13348 3556 13376
rect 3384 13336 3390 13348
rect 3528 13317 3556 13348
rect 1397 13311 1455 13317
rect 1397 13308 1409 13311
rect 900 13280 1409 13308
rect 900 13268 906 13280
rect 1397 13277 1409 13280
rect 1443 13277 1455 13311
rect 1397 13271 1455 13277
rect 2869 13311 2927 13317
rect 2869 13277 2881 13311
rect 2915 13277 2927 13311
rect 2869 13271 2927 13277
rect 3145 13311 3203 13317
rect 3145 13277 3157 13311
rect 3191 13308 3203 13311
rect 3421 13311 3479 13317
rect 3421 13308 3433 13311
rect 3191 13280 3433 13308
rect 3191 13277 3203 13280
rect 3145 13271 3203 13277
rect 3421 13277 3433 13280
rect 3467 13277 3479 13311
rect 3421 13271 3479 13277
rect 3513 13311 3571 13317
rect 3513 13277 3525 13311
rect 3559 13308 3571 13311
rect 3970 13308 3976 13320
rect 3559 13280 3976 13308
rect 3559 13277 3571 13280
rect 3513 13271 3571 13277
rect 2884 13240 2912 13271
rect 3970 13268 3976 13280
rect 4028 13268 4034 13320
rect 3234 13240 3240 13252
rect 2884 13212 3240 13240
rect 3234 13200 3240 13212
rect 3292 13200 3298 13252
rect 3344 13212 3556 13240
rect 2682 13132 2688 13184
rect 2740 13132 2746 13184
rect 3053 13175 3111 13181
rect 3053 13141 3065 13175
rect 3099 13172 3111 13175
rect 3344 13172 3372 13212
rect 3528 13184 3556 13212
rect 3099 13144 3372 13172
rect 3099 13141 3111 13144
rect 3053 13135 3111 13141
rect 3418 13132 3424 13184
rect 3476 13132 3482 13184
rect 3510 13132 3516 13184
rect 3568 13132 3574 13184
rect 4632 13172 4660 13416
rect 5092 13416 6745 13444
rect 4985 13311 5043 13317
rect 4985 13277 4997 13311
rect 5031 13308 5043 13311
rect 5092 13308 5120 13416
rect 5445 13379 5503 13385
rect 5445 13345 5457 13379
rect 5491 13376 5503 13379
rect 6089 13379 6147 13385
rect 6089 13376 6101 13379
rect 5491 13348 6101 13376
rect 5491 13345 5503 13348
rect 5445 13339 5503 13345
rect 6089 13345 6101 13348
rect 6135 13345 6147 13379
rect 6089 13339 6147 13345
rect 5031 13280 5120 13308
rect 5169 13311 5227 13317
rect 5031 13277 5043 13280
rect 4985 13271 5043 13277
rect 5169 13277 5181 13311
rect 5215 13308 5227 13311
rect 5460 13308 5488 13339
rect 5215 13280 5488 13308
rect 5215 13277 5227 13280
rect 5169 13271 5227 13277
rect 5534 13268 5540 13320
rect 5592 13268 5598 13320
rect 5905 13311 5963 13317
rect 5905 13277 5917 13311
rect 5951 13308 5963 13311
rect 6196 13308 6224 13416
rect 6733 13413 6745 13416
rect 6779 13413 6791 13447
rect 6733 13407 6791 13413
rect 8297 13447 8355 13453
rect 8297 13413 8309 13447
rect 8343 13413 8355 13447
rect 8297 13407 8355 13413
rect 8110 13376 8116 13388
rect 7852 13348 8116 13376
rect 5951 13280 6224 13308
rect 5951 13277 5963 13280
rect 5905 13271 5963 13277
rect 6270 13268 6276 13320
rect 6328 13268 6334 13320
rect 6362 13268 6368 13320
rect 6420 13308 6426 13320
rect 6549 13311 6607 13317
rect 6549 13308 6561 13311
rect 6420 13280 6561 13308
rect 6420 13268 6426 13280
rect 6549 13277 6561 13280
rect 6595 13308 6607 13311
rect 6825 13311 6883 13317
rect 6825 13308 6837 13311
rect 6595 13280 6837 13308
rect 6595 13277 6607 13280
rect 6549 13271 6607 13277
rect 6825 13277 6837 13280
rect 6871 13277 6883 13311
rect 6825 13271 6883 13277
rect 6914 13268 6920 13320
rect 6972 13308 6978 13320
rect 6972 13280 7328 13308
rect 6972 13268 6978 13280
rect 4706 13200 4712 13252
rect 4764 13240 4770 13252
rect 5261 13243 5319 13249
rect 5261 13240 5273 13243
rect 4764 13212 5273 13240
rect 4764 13200 4770 13212
rect 5261 13209 5273 13212
rect 5307 13209 5319 13243
rect 6288 13240 6316 13268
rect 6641 13243 6699 13249
rect 6641 13240 6653 13243
rect 6288 13212 6653 13240
rect 5261 13203 5319 13209
rect 6641 13209 6653 13212
rect 6687 13209 6699 13243
rect 7300 13240 7328 13280
rect 7374 13268 7380 13320
rect 7432 13308 7438 13320
rect 7852 13317 7880 13348
rect 8110 13336 8116 13348
rect 8168 13376 8174 13388
rect 8312 13376 8340 13407
rect 10410 13404 10416 13456
rect 10468 13444 10474 13456
rect 11333 13447 11391 13453
rect 11333 13444 11345 13447
rect 10468 13416 11345 13444
rect 10468 13404 10474 13416
rect 8570 13376 8576 13388
rect 8168 13348 8340 13376
rect 8404 13348 8576 13376
rect 8168 13336 8174 13348
rect 8404 13317 8432 13348
rect 8570 13336 8576 13348
rect 8628 13336 8634 13388
rect 10229 13379 10287 13385
rect 10229 13345 10241 13379
rect 10275 13376 10287 13379
rect 10318 13376 10324 13388
rect 10275 13348 10324 13376
rect 10275 13345 10287 13348
rect 10229 13339 10287 13345
rect 10318 13336 10324 13348
rect 10376 13336 10382 13388
rect 10612 13385 10640 13416
rect 11333 13413 11345 13416
rect 11379 13413 11391 13447
rect 11333 13407 11391 13413
rect 11606 13404 11612 13456
rect 11664 13444 11670 13456
rect 12618 13444 12624 13456
rect 11664 13416 12624 13444
rect 11664 13404 11670 13416
rect 12618 13404 12624 13416
rect 12676 13444 12682 13456
rect 12676 13416 13768 13444
rect 12676 13404 12682 13416
rect 10597 13379 10655 13385
rect 10597 13345 10609 13379
rect 10643 13345 10655 13379
rect 12434 13376 12440 13388
rect 10597 13339 10655 13345
rect 11072 13348 12440 13376
rect 11072 13320 11100 13348
rect 12434 13336 12440 13348
rect 12492 13336 12498 13388
rect 12912 13348 13676 13376
rect 7653 13311 7711 13317
rect 7653 13308 7665 13311
rect 7432 13280 7665 13308
rect 7432 13268 7438 13280
rect 7653 13277 7665 13280
rect 7699 13277 7711 13311
rect 7653 13271 7711 13277
rect 7837 13311 7895 13317
rect 7837 13277 7849 13311
rect 7883 13277 7895 13311
rect 7837 13271 7895 13277
rect 8297 13311 8355 13317
rect 8297 13277 8309 13311
rect 8343 13277 8355 13311
rect 8297 13271 8355 13277
rect 8389 13311 8447 13317
rect 8389 13277 8401 13311
rect 8435 13277 8447 13311
rect 8389 13271 8447 13277
rect 8496 13280 10088 13308
rect 8312 13240 8340 13271
rect 8496 13240 8524 13280
rect 7300 13212 8524 13240
rect 8573 13243 8631 13249
rect 6641 13203 6699 13209
rect 8573 13209 8585 13243
rect 8619 13240 8631 13243
rect 8938 13240 8944 13252
rect 8619 13212 8944 13240
rect 8619 13209 8631 13212
rect 8573 13203 8631 13209
rect 8938 13200 8944 13212
rect 8996 13200 9002 13252
rect 6362 13172 6368 13184
rect 4632 13144 6368 13172
rect 6362 13132 6368 13144
rect 6420 13132 6426 13184
rect 6454 13132 6460 13184
rect 6512 13132 6518 13184
rect 7558 13132 7564 13184
rect 7616 13172 7622 13184
rect 7653 13175 7711 13181
rect 7653 13172 7665 13175
rect 7616 13144 7665 13172
rect 7616 13132 7622 13144
rect 7653 13141 7665 13144
rect 7699 13141 7711 13175
rect 7653 13135 7711 13141
rect 9582 13132 9588 13184
rect 9640 13172 9646 13184
rect 9953 13175 10011 13181
rect 9953 13172 9965 13175
rect 9640 13144 9965 13172
rect 9640 13132 9646 13144
rect 9953 13141 9965 13144
rect 9999 13141 10011 13175
rect 10060 13172 10088 13280
rect 10134 13268 10140 13320
rect 10192 13308 10198 13320
rect 10689 13311 10747 13317
rect 10689 13308 10701 13311
rect 10192 13280 10701 13308
rect 10192 13268 10198 13280
rect 10689 13277 10701 13280
rect 10735 13277 10747 13311
rect 10689 13271 10747 13277
rect 10873 13311 10931 13317
rect 10873 13277 10885 13311
rect 10919 13277 10931 13311
rect 10873 13271 10931 13277
rect 10888 13240 10916 13271
rect 11054 13268 11060 13320
rect 11112 13268 11118 13320
rect 11149 13311 11207 13317
rect 11149 13277 11161 13311
rect 11195 13308 11207 13311
rect 11422 13308 11428 13320
rect 11195 13280 11428 13308
rect 11195 13277 11207 13280
rect 11149 13271 11207 13277
rect 11422 13268 11428 13280
rect 11480 13268 11486 13320
rect 11517 13311 11575 13317
rect 11517 13277 11529 13311
rect 11563 13308 11575 13311
rect 11606 13308 11612 13320
rect 11563 13280 11612 13308
rect 11563 13277 11575 13280
rect 11517 13271 11575 13277
rect 10962 13240 10968 13252
rect 10888 13212 10968 13240
rect 10962 13200 10968 13212
rect 11020 13240 11026 13252
rect 11241 13243 11299 13249
rect 11241 13240 11253 13243
rect 11020 13212 11253 13240
rect 11020 13200 11026 13212
rect 11241 13209 11253 13212
rect 11287 13209 11299 13243
rect 11241 13203 11299 13209
rect 11532 13172 11560 13271
rect 11606 13268 11612 13280
rect 11664 13268 11670 13320
rect 12452 13240 12480 13336
rect 12912 13317 12940 13348
rect 12897 13311 12955 13317
rect 12897 13277 12909 13311
rect 12943 13277 12955 13311
rect 12897 13271 12955 13277
rect 13170 13268 13176 13320
rect 13228 13268 13234 13320
rect 13357 13311 13415 13317
rect 13357 13277 13369 13311
rect 13403 13308 13415 13311
rect 13538 13308 13544 13320
rect 13403 13280 13544 13308
rect 13403 13277 13415 13280
rect 13357 13271 13415 13277
rect 13538 13268 13544 13280
rect 13596 13268 13602 13320
rect 12989 13243 13047 13249
rect 12989 13240 13001 13243
rect 12452 13212 13001 13240
rect 12989 13209 13001 13212
rect 13035 13209 13047 13243
rect 13188 13240 13216 13268
rect 13648 13249 13676 13348
rect 13740 13317 13768 13416
rect 13725 13311 13783 13317
rect 13725 13277 13737 13311
rect 13771 13277 13783 13311
rect 13725 13271 13783 13277
rect 17034 13268 17040 13320
rect 17092 13268 17098 13320
rect 13449 13243 13507 13249
rect 13449 13240 13461 13243
rect 13188 13212 13461 13240
rect 12989 13203 13047 13209
rect 13449 13209 13461 13212
rect 13495 13209 13507 13243
rect 13449 13203 13507 13209
rect 13633 13243 13691 13249
rect 13633 13209 13645 13243
rect 13679 13240 13691 13243
rect 13679 13212 16896 13240
rect 13679 13209 13691 13212
rect 13633 13203 13691 13209
rect 10060 13144 11560 13172
rect 9953 13135 10011 13141
rect 13722 13132 13728 13184
rect 13780 13132 13786 13184
rect 16868 13181 16896 13212
rect 16853 13175 16911 13181
rect 16853 13141 16865 13175
rect 16899 13141 16911 13175
rect 16853 13135 16911 13141
rect 1104 13082 17388 13104
rect 1104 13030 3645 13082
rect 3697 13030 3709 13082
rect 3761 13030 3773 13082
rect 3825 13030 3837 13082
rect 3889 13030 3901 13082
rect 3953 13030 7716 13082
rect 7768 13030 7780 13082
rect 7832 13030 7844 13082
rect 7896 13030 7908 13082
rect 7960 13030 7972 13082
rect 8024 13030 11787 13082
rect 11839 13030 11851 13082
rect 11903 13030 11915 13082
rect 11967 13030 11979 13082
rect 12031 13030 12043 13082
rect 12095 13030 15858 13082
rect 15910 13030 15922 13082
rect 15974 13030 15986 13082
rect 16038 13030 16050 13082
rect 16102 13030 16114 13082
rect 16166 13030 17388 13082
rect 1104 13008 17388 13030
rect 3145 12971 3203 12977
rect 2792 12940 3004 12968
rect 2792 12844 2820 12940
rect 2976 12900 3004 12940
rect 3145 12937 3157 12971
rect 3191 12968 3203 12971
rect 3234 12968 3240 12980
rect 3191 12940 3240 12968
rect 3191 12937 3203 12940
rect 3145 12931 3203 12937
rect 3234 12928 3240 12940
rect 3292 12928 3298 12980
rect 6181 12971 6239 12977
rect 4264 12940 4844 12968
rect 4264 12900 4292 12940
rect 2898 12872 4292 12900
rect 4706 12860 4712 12912
rect 4764 12860 4770 12912
rect 4816 12900 4844 12940
rect 6181 12937 6193 12971
rect 6227 12968 6239 12971
rect 6270 12968 6276 12980
rect 6227 12940 6276 12968
rect 6227 12937 6239 12940
rect 6181 12931 6239 12937
rect 6270 12928 6276 12940
rect 6328 12928 6334 12980
rect 8938 12928 8944 12980
rect 8996 12928 9002 12980
rect 10962 12928 10968 12980
rect 11020 12968 11026 12980
rect 11057 12971 11115 12977
rect 11057 12968 11069 12971
rect 11020 12940 11069 12968
rect 11020 12928 11026 12940
rect 11057 12937 11069 12940
rect 11103 12937 11115 12971
rect 11057 12931 11115 12937
rect 13170 12928 13176 12980
rect 13228 12968 13234 12980
rect 13265 12971 13323 12977
rect 13265 12968 13277 12971
rect 13228 12940 13277 12968
rect 13228 12928 13234 12940
rect 13265 12937 13277 12940
rect 13311 12937 13323 12971
rect 13265 12931 13323 12937
rect 13722 12928 13728 12980
rect 13780 12968 13786 12980
rect 14001 12971 14059 12977
rect 14001 12968 14013 12971
rect 13780 12940 14013 12968
rect 13780 12928 13786 12940
rect 14001 12937 14013 12940
rect 14047 12937 14059 12971
rect 14001 12931 14059 12937
rect 5166 12900 5172 12912
rect 4816 12872 5172 12900
rect 5166 12860 5172 12872
rect 5224 12860 5230 12912
rect 8478 12860 8484 12912
rect 8536 12860 8542 12912
rect 9582 12860 9588 12912
rect 9640 12860 9646 12912
rect 10870 12900 10876 12912
rect 10810 12872 10876 12900
rect 10870 12860 10876 12872
rect 10928 12860 10934 12912
rect 1394 12792 1400 12844
rect 1452 12792 1458 12844
rect 2774 12792 2780 12844
rect 2832 12792 2838 12844
rect 3421 12835 3479 12841
rect 3421 12832 3433 12835
rect 2884 12804 3433 12832
rect 2884 12776 2912 12804
rect 3421 12801 3433 12804
rect 3467 12801 3479 12835
rect 3421 12795 3479 12801
rect 12894 12792 12900 12844
rect 12952 12792 12958 12844
rect 13538 12792 13544 12844
rect 13596 12792 13602 12844
rect 14274 12792 14280 12844
rect 14332 12792 14338 12844
rect 15654 12792 15660 12844
rect 15712 12792 15718 12844
rect 1670 12724 1676 12776
rect 1728 12724 1734 12776
rect 2866 12724 2872 12776
rect 2924 12724 2930 12776
rect 3326 12724 3332 12776
rect 3384 12724 3390 12776
rect 4430 12724 4436 12776
rect 4488 12764 4494 12776
rect 5258 12764 5264 12776
rect 4488 12736 5264 12764
rect 4488 12724 4494 12736
rect 5258 12724 5264 12736
rect 5316 12724 5322 12776
rect 6178 12724 6184 12776
rect 6236 12764 6242 12776
rect 6822 12764 6828 12776
rect 6236 12736 6828 12764
rect 6236 12724 6242 12736
rect 6822 12724 6828 12736
rect 6880 12764 6886 12776
rect 7193 12767 7251 12773
rect 7193 12764 7205 12767
rect 6880 12736 7205 12764
rect 6880 12724 6886 12736
rect 7193 12733 7205 12736
rect 7239 12733 7251 12767
rect 7193 12727 7251 12733
rect 7466 12724 7472 12776
rect 7524 12724 7530 12776
rect 9306 12724 9312 12776
rect 9364 12724 9370 12776
rect 11514 12724 11520 12776
rect 11572 12724 11578 12776
rect 11793 12767 11851 12773
rect 11793 12733 11805 12767
rect 11839 12764 11851 12767
rect 13357 12767 13415 12773
rect 13357 12764 13369 12767
rect 11839 12736 13369 12764
rect 11839 12733 11851 12736
rect 11793 12727 11851 12733
rect 13357 12733 13369 12736
rect 13403 12733 13415 12767
rect 13357 12727 13415 12733
rect 13633 12767 13691 12773
rect 13633 12733 13645 12767
rect 13679 12764 13691 12767
rect 13814 12764 13820 12776
rect 13679 12736 13820 12764
rect 13679 12733 13691 12736
rect 13633 12727 13691 12733
rect 13814 12724 13820 12736
rect 13872 12724 13878 12776
rect 14550 12724 14556 12776
rect 14608 12724 14614 12776
rect 3789 12699 3847 12705
rect 3789 12665 3801 12699
rect 3835 12696 3847 12699
rect 4062 12696 4068 12708
rect 3835 12668 4068 12696
rect 3835 12665 3847 12668
rect 3789 12659 3847 12665
rect 4062 12656 4068 12668
rect 4120 12656 4126 12708
rect 16022 12588 16028 12640
rect 16080 12588 16086 12640
rect 1104 12538 17388 12560
rect 1104 12486 2985 12538
rect 3037 12486 3049 12538
rect 3101 12486 3113 12538
rect 3165 12486 3177 12538
rect 3229 12486 3241 12538
rect 3293 12486 7056 12538
rect 7108 12486 7120 12538
rect 7172 12486 7184 12538
rect 7236 12486 7248 12538
rect 7300 12486 7312 12538
rect 7364 12486 11127 12538
rect 11179 12486 11191 12538
rect 11243 12486 11255 12538
rect 11307 12486 11319 12538
rect 11371 12486 11383 12538
rect 11435 12486 15198 12538
rect 15250 12486 15262 12538
rect 15314 12486 15326 12538
rect 15378 12486 15390 12538
rect 15442 12486 15454 12538
rect 15506 12486 17388 12538
rect 1104 12464 17388 12486
rect 1670 12384 1676 12436
rect 1728 12424 1734 12436
rect 2041 12427 2099 12433
rect 2041 12424 2053 12427
rect 1728 12396 2053 12424
rect 1728 12384 1734 12396
rect 2041 12393 2053 12396
rect 2087 12393 2099 12427
rect 2041 12387 2099 12393
rect 2869 12427 2927 12433
rect 2869 12393 2881 12427
rect 2915 12424 2927 12427
rect 3326 12424 3332 12436
rect 2915 12396 3332 12424
rect 2915 12393 2927 12396
rect 2869 12387 2927 12393
rect 3326 12384 3332 12396
rect 3384 12384 3390 12436
rect 5534 12384 5540 12436
rect 5592 12384 5598 12436
rect 7466 12384 7472 12436
rect 7524 12384 7530 12436
rect 10870 12384 10876 12436
rect 10928 12424 10934 12436
rect 12894 12424 12900 12436
rect 10928 12396 12900 12424
rect 10928 12384 10934 12396
rect 12894 12384 12900 12396
rect 12952 12384 12958 12436
rect 14550 12384 14556 12436
rect 14608 12384 14614 12436
rect 16206 12384 16212 12436
rect 16264 12384 16270 12436
rect 8297 12359 8355 12365
rect 8297 12356 8309 12359
rect 7668 12328 8309 12356
rect 2225 12291 2283 12297
rect 2225 12257 2237 12291
rect 2271 12288 2283 12291
rect 2271 12260 2636 12288
rect 2271 12257 2283 12260
rect 2225 12251 2283 12257
rect 2317 12223 2375 12229
rect 2317 12189 2329 12223
rect 2363 12189 2375 12223
rect 2608 12220 2636 12260
rect 4062 12248 4068 12300
rect 4120 12248 4126 12300
rect 7374 12248 7380 12300
rect 7432 12288 7438 12300
rect 7668 12297 7696 12328
rect 8297 12325 8309 12328
rect 8343 12325 8355 12359
rect 8297 12319 8355 12325
rect 13357 12359 13415 12365
rect 13357 12325 13369 12359
rect 13403 12356 13415 12359
rect 13403 12328 14228 12356
rect 13403 12325 13415 12328
rect 13357 12319 13415 12325
rect 7653 12291 7711 12297
rect 7653 12288 7665 12291
rect 7432 12260 7665 12288
rect 7432 12248 7438 12260
rect 7653 12257 7665 12260
rect 7699 12257 7711 12291
rect 7653 12251 7711 12257
rect 8110 12248 8116 12300
rect 8168 12248 8174 12300
rect 8938 12288 8944 12300
rect 8496 12260 8944 12288
rect 2682 12220 2688 12232
rect 2608 12192 2688 12220
rect 2317 12183 2375 12189
rect 2332 12152 2360 12183
rect 2682 12180 2688 12192
rect 2740 12220 2746 12232
rect 2777 12223 2835 12229
rect 2777 12220 2789 12223
rect 2740 12192 2789 12220
rect 2740 12180 2746 12192
rect 2777 12189 2789 12192
rect 2823 12189 2835 12223
rect 2777 12183 2835 12189
rect 2961 12223 3019 12229
rect 2961 12189 2973 12223
rect 3007 12220 3019 12223
rect 3418 12220 3424 12232
rect 3007 12192 3424 12220
rect 3007 12189 3019 12192
rect 2961 12183 3019 12189
rect 2866 12152 2872 12164
rect 2332 12124 2872 12152
rect 2866 12112 2872 12124
rect 2924 12112 2930 12164
rect 2685 12087 2743 12093
rect 2685 12053 2697 12087
rect 2731 12084 2743 12087
rect 2976 12084 3004 12183
rect 3418 12180 3424 12192
rect 3476 12180 3482 12232
rect 3789 12223 3847 12229
rect 3789 12189 3801 12223
rect 3835 12189 3847 12223
rect 3789 12183 3847 12189
rect 3804 12152 3832 12183
rect 5166 12180 5172 12232
rect 5224 12180 5230 12232
rect 7745 12223 7803 12229
rect 7745 12189 7757 12223
rect 7791 12220 7803 12223
rect 8202 12220 8208 12232
rect 7791 12192 8208 12220
rect 7791 12189 7803 12192
rect 7745 12183 7803 12189
rect 8202 12180 8208 12192
rect 8260 12180 8266 12232
rect 8496 12229 8524 12260
rect 8938 12248 8944 12260
rect 8996 12248 9002 12300
rect 13538 12288 13544 12300
rect 13280 12260 13544 12288
rect 8481 12223 8539 12229
rect 8481 12189 8493 12223
rect 8527 12189 8539 12223
rect 8481 12183 8539 12189
rect 8662 12180 8668 12232
rect 8720 12220 8726 12232
rect 13280 12229 13308 12260
rect 13538 12248 13544 12260
rect 13596 12248 13602 12300
rect 14200 12297 14228 12328
rect 14185 12291 14243 12297
rect 14185 12257 14197 12291
rect 14231 12257 14243 12291
rect 14185 12251 14243 12257
rect 15841 12291 15899 12297
rect 15841 12257 15853 12291
rect 15887 12288 15899 12291
rect 16485 12291 16543 12297
rect 16485 12288 16497 12291
rect 15887 12260 16497 12288
rect 15887 12257 15899 12260
rect 15841 12251 15899 12257
rect 16485 12257 16497 12260
rect 16531 12257 16543 12291
rect 16485 12251 16543 12257
rect 8757 12223 8815 12229
rect 8757 12220 8769 12223
rect 8720 12192 8769 12220
rect 8720 12180 8726 12192
rect 8757 12189 8769 12192
rect 8803 12189 8815 12223
rect 8757 12183 8815 12189
rect 13265 12223 13323 12229
rect 13265 12189 13277 12223
rect 13311 12189 13323 12223
rect 13265 12183 13323 12189
rect 13449 12223 13507 12229
rect 13449 12189 13461 12223
rect 13495 12220 13507 12223
rect 13722 12220 13728 12232
rect 13495 12192 13728 12220
rect 13495 12189 13507 12192
rect 13449 12183 13507 12189
rect 13722 12180 13728 12192
rect 13780 12180 13786 12232
rect 13814 12180 13820 12232
rect 13872 12220 13878 12232
rect 14277 12223 14335 12229
rect 14277 12220 14289 12223
rect 13872 12192 14289 12220
rect 13872 12180 13878 12192
rect 14277 12189 14289 12192
rect 14323 12220 14335 12223
rect 15102 12220 15108 12232
rect 14323 12192 15108 12220
rect 14323 12189 14335 12192
rect 14277 12183 14335 12189
rect 15102 12180 15108 12192
rect 15160 12180 15166 12232
rect 15746 12180 15752 12232
rect 15804 12220 15810 12232
rect 15933 12223 15991 12229
rect 15933 12220 15945 12223
rect 15804 12192 15945 12220
rect 15804 12180 15810 12192
rect 15933 12189 15945 12192
rect 15979 12220 15991 12223
rect 16022 12220 16028 12232
rect 15979 12192 16028 12220
rect 15979 12189 15991 12192
rect 15933 12183 15991 12189
rect 16022 12180 16028 12192
rect 16080 12180 16086 12232
rect 16393 12223 16451 12229
rect 16393 12220 16405 12223
rect 16132 12192 16405 12220
rect 4338 12152 4344 12164
rect 3804 12124 4344 12152
rect 4338 12112 4344 12124
rect 4396 12112 4402 12164
rect 15562 12112 15568 12164
rect 15620 12152 15626 12164
rect 16132 12152 16160 12192
rect 16393 12189 16405 12192
rect 16439 12189 16451 12223
rect 16393 12183 16451 12189
rect 16577 12223 16635 12229
rect 16577 12189 16589 12223
rect 16623 12189 16635 12223
rect 16577 12183 16635 12189
rect 15620 12124 16160 12152
rect 15620 12112 15626 12124
rect 16206 12112 16212 12164
rect 16264 12152 16270 12164
rect 16592 12152 16620 12183
rect 16264 12124 16620 12152
rect 16264 12112 16270 12124
rect 2731 12056 3004 12084
rect 2731 12053 2743 12056
rect 2685 12047 2743 12053
rect 8662 12044 8668 12096
rect 8720 12044 8726 12096
rect 10226 12044 10232 12096
rect 10284 12084 10290 12096
rect 11054 12084 11060 12096
rect 10284 12056 11060 12084
rect 10284 12044 10290 12056
rect 11054 12044 11060 12056
rect 11112 12044 11118 12096
rect 1104 11994 17388 12016
rect 1104 11942 3645 11994
rect 3697 11942 3709 11994
rect 3761 11942 3773 11994
rect 3825 11942 3837 11994
rect 3889 11942 3901 11994
rect 3953 11942 7716 11994
rect 7768 11942 7780 11994
rect 7832 11942 7844 11994
rect 7896 11942 7908 11994
rect 7960 11942 7972 11994
rect 8024 11942 11787 11994
rect 11839 11942 11851 11994
rect 11903 11942 11915 11994
rect 11967 11942 11979 11994
rect 12031 11942 12043 11994
rect 12095 11942 15858 11994
rect 15910 11942 15922 11994
rect 15974 11942 15986 11994
rect 16038 11942 16050 11994
rect 16102 11942 16114 11994
rect 16166 11942 17388 11994
rect 1104 11920 17388 11942
rect 5994 11840 6000 11892
rect 6052 11880 6058 11892
rect 6454 11880 6460 11892
rect 6052 11852 6460 11880
rect 6052 11840 6058 11852
rect 6454 11840 6460 11852
rect 6512 11880 6518 11892
rect 8662 11880 8668 11892
rect 6512 11852 8668 11880
rect 6512 11840 6518 11852
rect 8662 11840 8668 11852
rect 8720 11880 8726 11892
rect 10226 11880 10232 11892
rect 8720 11852 10232 11880
rect 8720 11840 8726 11852
rect 10226 11840 10232 11852
rect 10284 11840 10290 11892
rect 10318 11840 10324 11892
rect 10376 11880 10382 11892
rect 10376 11852 14964 11880
rect 10376 11840 10382 11852
rect 9766 11772 9772 11824
rect 9824 11812 9830 11824
rect 13078 11812 13084 11824
rect 9824 11784 10640 11812
rect 13018 11784 13084 11812
rect 9824 11772 9830 11784
rect 4706 11704 4712 11756
rect 4764 11744 4770 11756
rect 4801 11747 4859 11753
rect 4801 11744 4813 11747
rect 4764 11716 4813 11744
rect 4764 11704 4770 11716
rect 4801 11713 4813 11716
rect 4847 11713 4859 11747
rect 4801 11707 4859 11713
rect 4985 11747 5043 11753
rect 4985 11713 4997 11747
rect 5031 11713 5043 11747
rect 4985 11707 5043 11713
rect 5721 11747 5779 11753
rect 5721 11713 5733 11747
rect 5767 11744 5779 11747
rect 5810 11744 5816 11756
rect 5767 11716 5816 11744
rect 5767 11713 5779 11716
rect 5721 11707 5779 11713
rect 5000 11676 5028 11707
rect 5810 11704 5816 11716
rect 5868 11704 5874 11756
rect 5902 11704 5908 11756
rect 5960 11704 5966 11756
rect 5997 11747 6055 11753
rect 5997 11713 6009 11747
rect 6043 11744 6055 11747
rect 6730 11744 6736 11756
rect 6043 11716 6736 11744
rect 6043 11713 6055 11716
rect 5997 11707 6055 11713
rect 6730 11704 6736 11716
rect 6788 11744 6794 11756
rect 6914 11744 6920 11756
rect 6788 11716 6920 11744
rect 6788 11704 6794 11716
rect 6914 11704 6920 11716
rect 6972 11704 6978 11756
rect 7469 11747 7527 11753
rect 7469 11713 7481 11747
rect 7515 11744 7527 11747
rect 8202 11744 8208 11756
rect 7515 11716 8208 11744
rect 7515 11713 7527 11716
rect 7469 11707 7527 11713
rect 8202 11704 8208 11716
rect 8260 11704 8266 11756
rect 10045 11747 10103 11753
rect 10045 11713 10057 11747
rect 10091 11713 10103 11747
rect 10045 11707 10103 11713
rect 5350 11676 5356 11688
rect 5000 11648 5356 11676
rect 5350 11636 5356 11648
rect 5408 11676 5414 11688
rect 5408 11648 5856 11676
rect 5408 11636 5414 11648
rect 5828 11617 5856 11648
rect 7558 11636 7564 11688
rect 7616 11636 7622 11688
rect 10060 11676 10088 11707
rect 10318 11704 10324 11756
rect 10376 11704 10382 11756
rect 10410 11704 10416 11756
rect 10468 11704 10474 11756
rect 10612 11753 10640 11784
rect 13078 11772 13084 11784
rect 13136 11812 13142 11824
rect 13722 11812 13728 11824
rect 13136 11784 13728 11812
rect 13136 11772 13142 11784
rect 13722 11772 13728 11784
rect 13780 11772 13786 11824
rect 14936 11812 14964 11852
rect 15102 11840 15108 11892
rect 15160 11840 15166 11892
rect 16301 11883 16359 11889
rect 16301 11880 16313 11883
rect 15212 11852 16313 11880
rect 15212 11812 15240 11852
rect 16301 11849 16313 11852
rect 16347 11849 16359 11883
rect 16301 11843 16359 11849
rect 14936 11784 15240 11812
rect 15746 11772 15752 11824
rect 15804 11812 15810 11824
rect 15804 11784 15884 11812
rect 15804 11772 15810 11784
rect 10597 11747 10655 11753
rect 10597 11713 10609 11747
rect 10643 11713 10655 11747
rect 10597 11707 10655 11713
rect 11514 11704 11520 11756
rect 11572 11704 11578 11756
rect 14918 11744 14924 11756
rect 14766 11730 14924 11744
rect 14752 11716 14924 11730
rect 10686 11676 10692 11688
rect 10060 11648 10692 11676
rect 10686 11636 10692 11648
rect 10744 11636 10750 11688
rect 11790 11636 11796 11688
rect 11848 11636 11854 11688
rect 13357 11679 13415 11685
rect 13357 11645 13369 11679
rect 13403 11645 13415 11679
rect 13357 11639 13415 11645
rect 5813 11611 5871 11617
rect 5813 11577 5825 11611
rect 5859 11577 5871 11611
rect 13372 11608 13400 11639
rect 13630 11636 13636 11688
rect 13688 11636 13694 11688
rect 13722 11636 13728 11688
rect 13780 11676 13786 11688
rect 14752 11676 14780 11716
rect 14918 11704 14924 11716
rect 14976 11704 14982 11756
rect 15856 11753 15884 11784
rect 15841 11747 15899 11753
rect 15841 11713 15853 11747
rect 15887 11713 15899 11747
rect 15841 11707 15899 11713
rect 16482 11704 16488 11756
rect 16540 11704 16546 11756
rect 16574 11704 16580 11756
rect 16632 11744 16638 11756
rect 16853 11747 16911 11753
rect 16853 11744 16865 11747
rect 16632 11716 16865 11744
rect 16632 11704 16638 11716
rect 16853 11713 16865 11716
rect 16899 11713 16911 11747
rect 16853 11707 16911 11713
rect 13780 11648 14780 11676
rect 13780 11636 13786 11648
rect 15562 11636 15568 11688
rect 15620 11676 15626 11688
rect 15749 11679 15807 11685
rect 15749 11676 15761 11679
rect 15620 11648 15761 11676
rect 15620 11636 15626 11648
rect 15749 11645 15761 11648
rect 15795 11645 15807 11679
rect 15749 11639 15807 11645
rect 16206 11636 16212 11688
rect 16264 11636 16270 11688
rect 5813 11571 5871 11577
rect 13188 11580 13400 11608
rect 4246 11500 4252 11552
rect 4304 11540 4310 11552
rect 4893 11543 4951 11549
rect 4893 11540 4905 11543
rect 4304 11512 4905 11540
rect 4304 11500 4310 11512
rect 4893 11509 4905 11512
rect 4939 11509 4951 11543
rect 4893 11503 4951 11509
rect 6914 11500 6920 11552
rect 6972 11540 6978 11552
rect 7193 11543 7251 11549
rect 7193 11540 7205 11543
rect 6972 11512 7205 11540
rect 6972 11500 6978 11512
rect 7193 11509 7205 11512
rect 7239 11509 7251 11543
rect 7193 11503 7251 11509
rect 9766 11500 9772 11552
rect 9824 11540 9830 11552
rect 9861 11543 9919 11549
rect 9861 11540 9873 11543
rect 9824 11512 9873 11540
rect 9824 11500 9830 11512
rect 9861 11509 9873 11512
rect 9907 11509 9919 11543
rect 9861 11503 9919 11509
rect 10505 11543 10563 11549
rect 10505 11509 10517 11543
rect 10551 11540 10563 11543
rect 10870 11540 10876 11552
rect 10551 11512 10876 11540
rect 10551 11509 10563 11512
rect 10505 11503 10563 11509
rect 10870 11500 10876 11512
rect 10928 11500 10934 11552
rect 11514 11500 11520 11552
rect 11572 11540 11578 11552
rect 13188 11540 13216 11580
rect 11572 11512 13216 11540
rect 11572 11500 11578 11512
rect 13262 11500 13268 11552
rect 13320 11500 13326 11552
rect 13372 11540 13400 11580
rect 15102 11540 15108 11552
rect 13372 11512 15108 11540
rect 15102 11500 15108 11512
rect 15160 11500 15166 11552
rect 15565 11543 15623 11549
rect 15565 11509 15577 11543
rect 15611 11540 15623 11543
rect 15654 11540 15660 11552
rect 15611 11512 15660 11540
rect 15611 11509 15623 11512
rect 15565 11503 15623 11509
rect 15654 11500 15660 11512
rect 15712 11500 15718 11552
rect 15746 11500 15752 11552
rect 15804 11540 15810 11552
rect 16761 11543 16819 11549
rect 16761 11540 16773 11543
rect 15804 11512 16773 11540
rect 15804 11500 15810 11512
rect 16761 11509 16773 11512
rect 16807 11509 16819 11543
rect 16761 11503 16819 11509
rect 1104 11450 17388 11472
rect 1104 11398 2985 11450
rect 3037 11398 3049 11450
rect 3101 11398 3113 11450
rect 3165 11398 3177 11450
rect 3229 11398 3241 11450
rect 3293 11398 7056 11450
rect 7108 11398 7120 11450
rect 7172 11398 7184 11450
rect 7236 11398 7248 11450
rect 7300 11398 7312 11450
rect 7364 11398 11127 11450
rect 11179 11398 11191 11450
rect 11243 11398 11255 11450
rect 11307 11398 11319 11450
rect 11371 11398 11383 11450
rect 11435 11398 15198 11450
rect 15250 11398 15262 11450
rect 15314 11398 15326 11450
rect 15378 11398 15390 11450
rect 15442 11398 15454 11450
rect 15506 11398 17388 11450
rect 1104 11376 17388 11398
rect 2866 11296 2872 11348
rect 2924 11336 2930 11348
rect 3145 11339 3203 11345
rect 3145 11336 3157 11339
rect 2924 11308 3157 11336
rect 2924 11296 2930 11308
rect 3145 11305 3157 11308
rect 3191 11305 3203 11339
rect 3145 11299 3203 11305
rect 5810 11296 5816 11348
rect 5868 11336 5874 11348
rect 6273 11339 6331 11345
rect 6273 11336 6285 11339
rect 5868 11308 6285 11336
rect 5868 11296 5874 11308
rect 6273 11305 6285 11308
rect 6319 11305 6331 11339
rect 6273 11299 6331 11305
rect 10686 11296 10692 11348
rect 10744 11296 10750 11348
rect 11241 11339 11299 11345
rect 11241 11305 11253 11339
rect 11287 11336 11299 11339
rect 11790 11336 11796 11348
rect 11287 11308 11796 11336
rect 11287 11305 11299 11308
rect 11241 11299 11299 11305
rect 11790 11296 11796 11308
rect 11848 11296 11854 11348
rect 12989 11339 13047 11345
rect 12989 11305 13001 11339
rect 13035 11336 13047 11339
rect 13630 11336 13636 11348
rect 13035 11308 13636 11336
rect 13035 11305 13047 11308
rect 12989 11299 13047 11305
rect 13630 11296 13636 11308
rect 13688 11296 13694 11348
rect 3789 11271 3847 11277
rect 3789 11268 3801 11271
rect 2746 11240 3801 11268
rect 1394 11160 1400 11212
rect 1452 11160 1458 11212
rect 1673 11203 1731 11209
rect 1673 11169 1685 11203
rect 1719 11200 1731 11203
rect 2746 11200 2774 11240
rect 3789 11237 3801 11240
rect 3835 11237 3847 11271
rect 3789 11231 3847 11237
rect 6914 11228 6920 11280
rect 6972 11228 6978 11280
rect 1719 11172 2774 11200
rect 1719 11169 1731 11172
rect 1673 11163 1731 11169
rect 4246 11160 4252 11212
rect 4304 11160 4310 11212
rect 4338 11160 4344 11212
rect 4396 11200 4402 11212
rect 4525 11203 4583 11209
rect 4525 11200 4537 11203
rect 4396 11172 4537 11200
rect 4396 11160 4402 11172
rect 4525 11169 4537 11172
rect 4571 11169 4583 11203
rect 4525 11163 4583 11169
rect 5166 11160 5172 11212
rect 5224 11200 5230 11212
rect 6932 11200 6960 11228
rect 7193 11203 7251 11209
rect 7193 11200 7205 11203
rect 5224 11172 6040 11200
rect 6932 11172 7205 11200
rect 5224 11160 5230 11172
rect 2774 11092 2780 11144
rect 2832 11092 2838 11144
rect 4154 11092 4160 11144
rect 4212 11092 4218 11144
rect 4798 11024 4804 11076
rect 4856 11024 4862 11076
rect 6012 11064 6040 11172
rect 7193 11169 7205 11172
rect 7239 11169 7251 11203
rect 8386 11200 8392 11212
rect 7193 11163 7251 11169
rect 8312 11172 8392 11200
rect 6822 11092 6828 11144
rect 6880 11132 6886 11144
rect 6917 11135 6975 11141
rect 6917 11132 6929 11135
rect 6880 11104 6929 11132
rect 6880 11092 6886 11104
rect 6917 11101 6929 11104
rect 6963 11101 6975 11135
rect 8312 11118 8340 11172
rect 8386 11160 8392 11172
rect 8444 11160 8450 11212
rect 8662 11160 8668 11212
rect 8720 11160 8726 11212
rect 8941 11203 8999 11209
rect 8941 11169 8953 11203
rect 8987 11200 8999 11203
rect 9306 11200 9312 11212
rect 8987 11172 9312 11200
rect 8987 11169 8999 11172
rect 8941 11163 8999 11169
rect 9306 11160 9312 11172
rect 9364 11160 9370 11212
rect 10870 11160 10876 11212
rect 10928 11160 10934 11212
rect 12802 11160 12808 11212
rect 12860 11160 12866 11212
rect 14274 11160 14280 11212
rect 14332 11200 14338 11212
rect 15013 11203 15071 11209
rect 15013 11200 15025 11203
rect 14332 11172 15025 11200
rect 14332 11160 14338 11172
rect 15013 11169 15025 11172
rect 15059 11169 15071 11203
rect 15013 11163 15071 11169
rect 15289 11203 15347 11209
rect 15289 11169 15301 11203
rect 15335 11200 15347 11203
rect 15654 11200 15660 11212
rect 15335 11172 15660 11200
rect 15335 11169 15347 11172
rect 15289 11163 15347 11169
rect 15654 11160 15660 11172
rect 15712 11160 15718 11212
rect 16482 11160 16488 11212
rect 16540 11200 16546 11212
rect 16761 11203 16819 11209
rect 16761 11200 16773 11203
rect 16540 11172 16773 11200
rect 16540 11160 16546 11172
rect 16761 11169 16773 11172
rect 16807 11169 16819 11203
rect 16761 11163 16819 11169
rect 6917 11095 6975 11101
rect 10962 11092 10968 11144
rect 11020 11092 11026 11144
rect 12434 11092 12440 11144
rect 12492 11132 12498 11144
rect 12713 11135 12771 11141
rect 12713 11132 12725 11135
rect 12492 11104 12725 11132
rect 12492 11092 12498 11104
rect 12713 11101 12725 11104
rect 12759 11132 12771 11135
rect 13262 11132 13268 11144
rect 12759 11104 13268 11132
rect 12759 11101 12771 11104
rect 12713 11095 12771 11101
rect 13262 11092 13268 11104
rect 13320 11092 13326 11144
rect 17034 11092 17040 11144
rect 17092 11092 17098 11144
rect 6365 11067 6423 11073
rect 6365 11064 6377 11067
rect 6012 11050 6377 11064
rect 6026 11036 6377 11050
rect 6365 11033 6377 11036
rect 6411 11033 6423 11067
rect 6365 11027 6423 11033
rect 6733 11067 6791 11073
rect 6733 11033 6745 11067
rect 6779 11064 6791 11067
rect 6779 11036 7604 11064
rect 6779 11033 6791 11036
rect 6733 11027 6791 11033
rect 1394 10956 1400 11008
rect 1452 10996 1458 11008
rect 2590 10996 2596 11008
rect 1452 10968 2596 10996
rect 1452 10956 1458 10968
rect 2590 10956 2596 10968
rect 2648 10956 2654 11008
rect 7576 10996 7604 11036
rect 9214 11024 9220 11076
rect 9272 11024 9278 11076
rect 10778 11064 10784 11076
rect 10442 11036 10784 11064
rect 10778 11024 10784 11036
rect 10836 11024 10842 11076
rect 15746 11024 15752 11076
rect 15804 11024 15810 11076
rect 8478 10996 8484 11008
rect 7576 10968 8484 10996
rect 8478 10956 8484 10968
rect 8536 10996 8542 11008
rect 16574 10996 16580 11008
rect 8536 10968 16580 10996
rect 8536 10956 8542 10968
rect 16574 10956 16580 10968
rect 16632 10956 16638 11008
rect 16850 10956 16856 11008
rect 16908 10956 16914 11008
rect 1104 10906 17388 10928
rect 1104 10854 3645 10906
rect 3697 10854 3709 10906
rect 3761 10854 3773 10906
rect 3825 10854 3837 10906
rect 3889 10854 3901 10906
rect 3953 10854 7716 10906
rect 7768 10854 7780 10906
rect 7832 10854 7844 10906
rect 7896 10854 7908 10906
rect 7960 10854 7972 10906
rect 8024 10854 11787 10906
rect 11839 10854 11851 10906
rect 11903 10854 11915 10906
rect 11967 10854 11979 10906
rect 12031 10854 12043 10906
rect 12095 10854 15858 10906
rect 15910 10854 15922 10906
rect 15974 10854 15986 10906
rect 16038 10854 16050 10906
rect 16102 10854 16114 10906
rect 16166 10854 17388 10906
rect 1104 10832 17388 10854
rect 1581 10795 1639 10801
rect 1581 10761 1593 10795
rect 1627 10761 1639 10795
rect 1581 10755 1639 10761
rect 2501 10795 2559 10801
rect 2501 10761 2513 10795
rect 2547 10761 2559 10795
rect 2501 10755 2559 10761
rect 1596 10724 1624 10755
rect 2516 10724 2544 10755
rect 2774 10752 2780 10804
rect 2832 10792 2838 10804
rect 2832 10764 3280 10792
rect 2832 10752 2838 10764
rect 2869 10727 2927 10733
rect 2869 10724 2881 10727
rect 1596 10696 2360 10724
rect 2516 10696 2881 10724
rect 842 10616 848 10668
rect 900 10656 906 10668
rect 1397 10659 1455 10665
rect 1397 10656 1409 10659
rect 900 10628 1409 10656
rect 900 10616 906 10628
rect 1397 10625 1409 10628
rect 1443 10625 1455 10659
rect 1397 10619 1455 10625
rect 2038 10616 2044 10668
rect 2096 10656 2102 10668
rect 2133 10659 2191 10665
rect 2133 10656 2145 10659
rect 2096 10628 2145 10656
rect 2096 10616 2102 10628
rect 2133 10625 2145 10628
rect 2179 10625 2191 10659
rect 2133 10619 2191 10625
rect 2225 10591 2283 10597
rect 2225 10557 2237 10591
rect 2271 10557 2283 10591
rect 2225 10551 2283 10557
rect 2240 10452 2268 10551
rect 2332 10520 2360 10696
rect 2869 10693 2881 10696
rect 2915 10693 2927 10727
rect 3252 10724 3280 10764
rect 4154 10752 4160 10804
rect 4212 10792 4218 10804
rect 4341 10795 4399 10801
rect 4341 10792 4353 10795
rect 4212 10764 4353 10792
rect 4212 10752 4218 10764
rect 4341 10761 4353 10764
rect 4387 10761 4399 10795
rect 4341 10755 4399 10761
rect 4617 10795 4675 10801
rect 4617 10761 4629 10795
rect 4663 10792 4675 10795
rect 4798 10792 4804 10804
rect 4663 10764 4804 10792
rect 4663 10761 4675 10764
rect 4617 10755 4675 10761
rect 3252 10696 3358 10724
rect 2869 10687 2927 10693
rect 2590 10616 2596 10668
rect 2648 10616 2654 10668
rect 4356 10656 4384 10755
rect 4798 10752 4804 10764
rect 4856 10752 4862 10804
rect 5261 10795 5319 10801
rect 5261 10761 5273 10795
rect 5307 10792 5319 10795
rect 5350 10792 5356 10804
rect 5307 10764 5356 10792
rect 5307 10761 5319 10764
rect 5261 10755 5319 10761
rect 5350 10752 5356 10764
rect 5408 10752 5414 10804
rect 6730 10752 6736 10804
rect 6788 10792 6794 10804
rect 7929 10795 7987 10801
rect 7929 10792 7941 10795
rect 6788 10764 7941 10792
rect 6788 10752 6794 10764
rect 7929 10761 7941 10764
rect 7975 10761 7987 10795
rect 7929 10755 7987 10761
rect 8205 10795 8263 10801
rect 8205 10761 8217 10795
rect 8251 10792 8263 10795
rect 8386 10792 8392 10804
rect 8251 10764 8392 10792
rect 8251 10761 8263 10764
rect 8205 10755 8263 10761
rect 5997 10727 6055 10733
rect 5997 10693 6009 10727
rect 6043 10724 6055 10727
rect 6043 10696 7328 10724
rect 6043 10693 6055 10696
rect 5997 10687 6055 10693
rect 4893 10659 4951 10665
rect 4893 10656 4905 10659
rect 4356 10628 4905 10656
rect 4893 10625 4905 10628
rect 4939 10625 4951 10659
rect 4893 10619 4951 10625
rect 5810 10616 5816 10668
rect 5868 10616 5874 10668
rect 7300 10665 7328 10696
rect 6089 10659 6147 10665
rect 6089 10625 6101 10659
rect 6135 10625 6147 10659
rect 6089 10619 6147 10625
rect 7285 10659 7343 10665
rect 7285 10625 7297 10659
rect 7331 10656 7343 10659
rect 7558 10656 7564 10668
rect 7331 10628 7564 10656
rect 7331 10625 7343 10628
rect 7285 10619 7343 10625
rect 2700 10560 4660 10588
rect 2700 10520 2728 10560
rect 2332 10492 2728 10520
rect 4632 10520 4660 10560
rect 4706 10548 4712 10600
rect 4764 10588 4770 10600
rect 4801 10591 4859 10597
rect 4801 10588 4813 10591
rect 4764 10560 4813 10588
rect 4764 10548 4770 10560
rect 4801 10557 4813 10560
rect 4847 10588 4859 10591
rect 5629 10591 5687 10597
rect 5629 10588 5641 10591
rect 4847 10560 5641 10588
rect 4847 10557 4859 10560
rect 4801 10551 4859 10557
rect 5629 10557 5641 10560
rect 5675 10557 5687 10591
rect 5629 10551 5687 10557
rect 5902 10520 5908 10532
rect 4632 10492 5908 10520
rect 5902 10480 5908 10492
rect 5960 10520 5966 10532
rect 6104 10520 6132 10619
rect 7558 10616 7564 10628
rect 7616 10656 7622 10668
rect 7745 10659 7803 10665
rect 7745 10656 7757 10659
rect 7616 10628 7757 10656
rect 7616 10616 7622 10628
rect 7745 10625 7757 10628
rect 7791 10625 7803 10659
rect 7944 10656 7972 10755
rect 8386 10752 8392 10764
rect 8444 10752 8450 10804
rect 9214 10752 9220 10804
rect 9272 10792 9278 10804
rect 9585 10795 9643 10801
rect 9585 10792 9597 10795
rect 9272 10764 9597 10792
rect 9272 10752 9278 10764
rect 9585 10761 9597 10764
rect 9631 10761 9643 10795
rect 9585 10755 9643 10761
rect 10229 10795 10287 10801
rect 10229 10761 10241 10795
rect 10275 10792 10287 10795
rect 10410 10792 10416 10804
rect 10275 10764 10416 10792
rect 10275 10761 10287 10764
rect 10229 10755 10287 10761
rect 10410 10752 10416 10764
rect 10468 10752 10474 10804
rect 12802 10752 12808 10804
rect 12860 10792 12866 10804
rect 12989 10795 13047 10801
rect 12989 10792 13001 10795
rect 12860 10764 13001 10792
rect 12860 10752 12866 10764
rect 12989 10761 13001 10764
rect 13035 10761 13047 10795
rect 12989 10755 13047 10761
rect 14918 10752 14924 10804
rect 14976 10792 14982 10804
rect 15749 10795 15807 10801
rect 15749 10792 15761 10795
rect 14976 10764 15761 10792
rect 14976 10752 14982 10764
rect 15749 10761 15761 10764
rect 15795 10761 15807 10795
rect 15749 10755 15807 10761
rect 16206 10752 16212 10804
rect 16264 10752 16270 10804
rect 16574 10792 16580 10804
rect 16316 10764 16580 10792
rect 8297 10727 8355 10733
rect 8297 10693 8309 10727
rect 8343 10724 8355 10727
rect 8478 10724 8484 10736
rect 8343 10696 8484 10724
rect 8343 10693 8355 10696
rect 8297 10687 8355 10693
rect 8478 10684 8484 10696
rect 8536 10684 8542 10736
rect 10597 10727 10655 10733
rect 8772 10696 10364 10724
rect 8772 10668 8800 10696
rect 8754 10656 8760 10668
rect 7944 10628 8760 10656
rect 7745 10619 7803 10625
rect 8754 10616 8760 10628
rect 8812 10616 8818 10668
rect 9766 10616 9772 10668
rect 9824 10616 9830 10668
rect 10336 10665 10364 10696
rect 10597 10693 10609 10727
rect 10643 10724 10655 10727
rect 10686 10724 10692 10736
rect 10643 10696 10692 10724
rect 10643 10693 10655 10696
rect 10597 10687 10655 10693
rect 10686 10684 10692 10696
rect 10744 10684 10750 10736
rect 14936 10724 14964 10752
rect 12360 10696 13124 10724
rect 14858 10696 14964 10724
rect 10321 10659 10379 10665
rect 10321 10625 10333 10659
rect 10367 10625 10379 10659
rect 10321 10619 10379 10625
rect 10410 10616 10416 10668
rect 10468 10616 10474 10668
rect 12360 10665 12388 10696
rect 12345 10659 12403 10665
rect 12345 10625 12357 10659
rect 12391 10625 12403 10659
rect 12345 10619 12403 10625
rect 12434 10616 12440 10668
rect 12492 10616 12498 10668
rect 13096 10665 13124 10696
rect 15194 10684 15200 10736
rect 15252 10724 15258 10736
rect 16025 10727 16083 10733
rect 15252 10696 15608 10724
rect 15252 10684 15258 10696
rect 12897 10659 12955 10665
rect 12897 10656 12909 10659
rect 12820 10628 12909 10656
rect 12820 10600 12848 10628
rect 12897 10625 12909 10628
rect 12943 10625 12955 10659
rect 12897 10619 12955 10625
rect 13081 10659 13139 10665
rect 13081 10625 13093 10659
rect 13127 10656 13139 10659
rect 13262 10656 13268 10668
rect 13127 10628 13268 10656
rect 13127 10625 13139 10628
rect 13081 10619 13139 10625
rect 13262 10616 13268 10628
rect 13320 10616 13326 10668
rect 15580 10665 15608 10696
rect 16025 10693 16037 10727
rect 16071 10724 16083 10727
rect 16316 10724 16344 10764
rect 16574 10752 16580 10764
rect 16632 10752 16638 10804
rect 16071 10696 16344 10724
rect 16071 10693 16083 10696
rect 16025 10687 16083 10693
rect 16482 10684 16488 10736
rect 16540 10684 16546 10736
rect 15565 10659 15623 10665
rect 15565 10625 15577 10659
rect 15611 10625 15623 10659
rect 15565 10619 15623 10625
rect 16209 10659 16267 10665
rect 16209 10625 16221 10659
rect 16255 10625 16267 10659
rect 16209 10619 16267 10625
rect 16301 10659 16359 10665
rect 16301 10625 16313 10659
rect 16347 10656 16359 10659
rect 16850 10656 16856 10668
rect 16347 10628 16856 10656
rect 16347 10625 16359 10628
rect 16301 10619 16359 10625
rect 9861 10591 9919 10597
rect 9861 10557 9873 10591
rect 9907 10557 9919 10591
rect 9861 10551 9919 10557
rect 5960 10492 6132 10520
rect 9876 10520 9904 10551
rect 12802 10548 12808 10600
rect 12860 10548 12866 10600
rect 14918 10548 14924 10600
rect 14976 10588 14982 10600
rect 15289 10591 15347 10597
rect 15289 10588 15301 10591
rect 14976 10560 15301 10588
rect 14976 10548 14982 10560
rect 15289 10557 15301 10560
rect 15335 10557 15347 10591
rect 16224 10588 16252 10619
rect 16850 10616 16856 10628
rect 16908 10616 16914 10668
rect 17034 10616 17040 10668
rect 17092 10616 17098 10668
rect 16942 10588 16948 10600
rect 16224 10560 16948 10588
rect 15289 10551 15347 10557
rect 16942 10548 16948 10560
rect 17000 10548 17006 10600
rect 10962 10520 10968 10532
rect 9876 10492 10968 10520
rect 5960 10480 5966 10492
rect 10962 10480 10968 10492
rect 11020 10520 11026 10532
rect 13817 10523 13875 10529
rect 13817 10520 13829 10523
rect 11020 10492 13829 10520
rect 11020 10480 11026 10492
rect 13817 10489 13829 10492
rect 13863 10489 13875 10523
rect 16853 10523 16911 10529
rect 16853 10520 16865 10523
rect 13817 10483 13875 10489
rect 15488 10492 16865 10520
rect 2866 10452 2872 10464
rect 2240 10424 2872 10452
rect 2866 10412 2872 10424
rect 2924 10412 2930 10464
rect 7561 10455 7619 10461
rect 7561 10421 7573 10455
rect 7607 10452 7619 10455
rect 8202 10452 8208 10464
rect 7607 10424 8208 10452
rect 7607 10421 7619 10424
rect 7561 10415 7619 10421
rect 8202 10412 8208 10424
rect 8260 10412 8266 10464
rect 11698 10412 11704 10464
rect 11756 10452 11762 10464
rect 12161 10455 12219 10461
rect 12161 10452 12173 10455
rect 11756 10424 12173 10452
rect 11756 10412 11762 10424
rect 12161 10421 12173 10424
rect 12207 10421 12219 10455
rect 12161 10415 12219 10421
rect 13722 10412 13728 10464
rect 13780 10452 13786 10464
rect 15488 10452 15516 10492
rect 16853 10489 16865 10492
rect 16899 10489 16911 10523
rect 16853 10483 16911 10489
rect 13780 10424 15516 10452
rect 13780 10412 13786 10424
rect 1104 10362 17388 10384
rect 1104 10310 2985 10362
rect 3037 10310 3049 10362
rect 3101 10310 3113 10362
rect 3165 10310 3177 10362
rect 3229 10310 3241 10362
rect 3293 10310 7056 10362
rect 7108 10310 7120 10362
rect 7172 10310 7184 10362
rect 7236 10310 7248 10362
rect 7300 10310 7312 10362
rect 7364 10310 11127 10362
rect 11179 10310 11191 10362
rect 11243 10310 11255 10362
rect 11307 10310 11319 10362
rect 11371 10310 11383 10362
rect 11435 10310 15198 10362
rect 15250 10310 15262 10362
rect 15314 10310 15326 10362
rect 15378 10310 15390 10362
rect 15442 10310 15454 10362
rect 15506 10310 17388 10362
rect 1104 10288 17388 10310
rect 13262 10208 13268 10260
rect 13320 10208 13326 10260
rect 14918 10208 14924 10260
rect 14976 10248 14982 10260
rect 15013 10251 15071 10257
rect 15013 10248 15025 10251
rect 14976 10220 15025 10248
rect 14976 10208 14982 10220
rect 15013 10217 15025 10220
rect 15059 10217 15071 10251
rect 15013 10211 15071 10217
rect 15562 10208 15568 10260
rect 15620 10248 15626 10260
rect 16117 10251 16175 10257
rect 16117 10248 16129 10251
rect 15620 10220 16129 10248
rect 15620 10208 15626 10220
rect 16117 10217 16129 10220
rect 16163 10217 16175 10251
rect 16117 10211 16175 10217
rect 11698 10072 11704 10124
rect 11756 10072 11762 10124
rect 13078 10072 13084 10124
rect 13136 10112 13142 10124
rect 13173 10115 13231 10121
rect 13173 10112 13185 10115
rect 13136 10084 13185 10112
rect 13136 10072 13142 10084
rect 13173 10081 13185 10084
rect 13219 10112 13231 10115
rect 13219 10084 13492 10112
rect 13219 10081 13231 10084
rect 13173 10075 13231 10081
rect 1394 10004 1400 10056
rect 1452 10004 1458 10056
rect 8021 10047 8079 10053
rect 8021 10013 8033 10047
rect 8067 10044 8079 10047
rect 8110 10044 8116 10056
rect 8067 10016 8116 10044
rect 8067 10013 8079 10016
rect 8021 10007 8079 10013
rect 8110 10004 8116 10016
rect 8168 10004 8174 10056
rect 8205 10047 8263 10053
rect 8205 10013 8217 10047
rect 8251 10044 8263 10047
rect 8294 10044 8300 10056
rect 8251 10016 8300 10044
rect 8251 10013 8263 10016
rect 8205 10007 8263 10013
rect 8294 10004 8300 10016
rect 8352 10004 8358 10056
rect 11422 10004 11428 10056
rect 11480 10004 11486 10056
rect 13464 10053 13492 10084
rect 15378 10072 15384 10124
rect 15436 10072 15442 10124
rect 13449 10047 13507 10053
rect 13449 10013 13461 10047
rect 13495 10013 13507 10047
rect 13449 10007 13507 10013
rect 13722 10004 13728 10056
rect 13780 10004 13786 10056
rect 15289 10047 15347 10053
rect 15289 10013 15301 10047
rect 15335 10044 15347 10047
rect 15746 10044 15752 10056
rect 15335 10016 15752 10044
rect 15335 10013 15347 10016
rect 15289 10007 15347 10013
rect 15746 10004 15752 10016
rect 15804 10004 15810 10056
rect 16301 10047 16359 10053
rect 16301 10013 16313 10047
rect 16347 10044 16359 10047
rect 16482 10044 16488 10056
rect 16347 10016 16488 10044
rect 16347 10013 16359 10016
rect 16301 10007 16359 10013
rect 16482 10004 16488 10016
rect 16540 10004 16546 10056
rect 16577 10047 16635 10053
rect 16577 10013 16589 10047
rect 16623 10044 16635 10047
rect 16850 10044 16856 10056
rect 16623 10016 16856 10044
rect 16623 10013 16635 10016
rect 16577 10007 16635 10013
rect 16850 10004 16856 10016
rect 16908 10004 16914 10056
rect 12434 9936 12440 9988
rect 12492 9936 12498 9988
rect 1581 9911 1639 9917
rect 1581 9877 1593 9911
rect 1627 9908 1639 9911
rect 2958 9908 2964 9920
rect 1627 9880 2964 9908
rect 1627 9877 1639 9880
rect 1581 9871 1639 9877
rect 2958 9868 2964 9880
rect 3016 9868 3022 9920
rect 8113 9911 8171 9917
rect 8113 9877 8125 9911
rect 8159 9908 8171 9911
rect 8478 9908 8484 9920
rect 8159 9880 8484 9908
rect 8159 9877 8171 9880
rect 8113 9871 8171 9877
rect 8478 9868 8484 9880
rect 8536 9868 8542 9920
rect 12710 9868 12716 9920
rect 12768 9908 12774 9920
rect 13633 9911 13691 9917
rect 13633 9908 13645 9911
rect 12768 9880 13645 9908
rect 12768 9868 12774 9880
rect 13633 9877 13645 9880
rect 13679 9877 13691 9911
rect 13633 9871 13691 9877
rect 16206 9868 16212 9920
rect 16264 9908 16270 9920
rect 16485 9911 16543 9917
rect 16485 9908 16497 9911
rect 16264 9880 16497 9908
rect 16264 9868 16270 9880
rect 16485 9877 16497 9880
rect 16531 9877 16543 9911
rect 16485 9871 16543 9877
rect 1104 9818 17388 9840
rect 1104 9766 3645 9818
rect 3697 9766 3709 9818
rect 3761 9766 3773 9818
rect 3825 9766 3837 9818
rect 3889 9766 3901 9818
rect 3953 9766 7716 9818
rect 7768 9766 7780 9818
rect 7832 9766 7844 9818
rect 7896 9766 7908 9818
rect 7960 9766 7972 9818
rect 8024 9766 11787 9818
rect 11839 9766 11851 9818
rect 11903 9766 11915 9818
rect 11967 9766 11979 9818
rect 12031 9766 12043 9818
rect 12095 9766 15858 9818
rect 15910 9766 15922 9818
rect 15974 9766 15986 9818
rect 16038 9766 16050 9818
rect 16102 9766 16114 9818
rect 16166 9766 17388 9818
rect 1104 9744 17388 9766
rect 2866 9664 2872 9716
rect 2924 9704 2930 9716
rect 3053 9707 3111 9713
rect 3053 9704 3065 9707
rect 2924 9676 3065 9704
rect 2924 9664 2930 9676
rect 3053 9673 3065 9676
rect 3099 9673 3111 9707
rect 3053 9667 3111 9673
rect 12802 9664 12808 9716
rect 12860 9664 12866 9716
rect 15378 9664 15384 9716
rect 15436 9704 15442 9716
rect 15565 9707 15623 9713
rect 15565 9704 15577 9707
rect 15436 9676 15577 9704
rect 15436 9664 15442 9676
rect 15565 9673 15577 9676
rect 15611 9673 15623 9707
rect 15565 9667 15623 9673
rect 16206 9664 16212 9716
rect 16264 9704 16270 9716
rect 16393 9707 16451 9713
rect 16393 9704 16405 9707
rect 16264 9676 16405 9704
rect 16264 9664 16270 9676
rect 16393 9673 16405 9676
rect 16439 9673 16451 9707
rect 16393 9667 16451 9673
rect 1578 9596 1584 9648
rect 1636 9596 1642 9648
rect 3510 9596 3516 9648
rect 3568 9636 3574 9648
rect 3970 9636 3976 9648
rect 3568 9608 3976 9636
rect 3568 9596 3574 9608
rect 3970 9596 3976 9608
rect 4028 9636 4034 9648
rect 8202 9636 8208 9648
rect 4028 9608 8208 9636
rect 4028 9596 4034 9608
rect 8202 9596 8208 9608
rect 8260 9596 8266 9648
rect 9950 9596 9956 9648
rect 10008 9596 10014 9648
rect 13078 9596 13084 9648
rect 13136 9596 13142 9648
rect 1949 9571 2007 9577
rect 1949 9537 1961 9571
rect 1995 9568 2007 9571
rect 1995 9540 2544 9568
rect 1995 9537 2007 9540
rect 1949 9531 2007 9537
rect 2038 9460 2044 9512
rect 2096 9460 2102 9512
rect 2406 9460 2412 9512
rect 2464 9460 2470 9512
rect 2516 9509 2544 9540
rect 2682 9528 2688 9580
rect 2740 9528 2746 9580
rect 2866 9528 2872 9580
rect 2924 9528 2930 9580
rect 2958 9528 2964 9580
rect 3016 9528 3022 9580
rect 3053 9571 3111 9577
rect 3053 9537 3065 9571
rect 3099 9566 3111 9571
rect 3237 9571 3295 9577
rect 3099 9538 3188 9566
rect 3099 9537 3111 9538
rect 3053 9531 3111 9537
rect 2501 9503 2559 9509
rect 2501 9469 2513 9503
rect 2547 9500 2559 9503
rect 2547 9472 2912 9500
rect 2547 9469 2559 9472
rect 2501 9463 2559 9469
rect 1578 9392 1584 9444
rect 1636 9432 1642 9444
rect 2884 9432 2912 9472
rect 3160 9432 3188 9538
rect 3237 9537 3249 9571
rect 3283 9568 3295 9571
rect 3326 9568 3332 9580
rect 3283 9540 3332 9568
rect 3283 9537 3295 9540
rect 3237 9531 3295 9537
rect 3326 9528 3332 9540
rect 3384 9528 3390 9580
rect 5718 9528 5724 9580
rect 5776 9528 5782 9580
rect 5810 9528 5816 9580
rect 5868 9528 5874 9580
rect 5997 9571 6055 9577
rect 5997 9537 6009 9571
rect 6043 9537 6055 9571
rect 5997 9531 6055 9537
rect 7837 9571 7895 9577
rect 7837 9537 7849 9571
rect 7883 9568 7895 9571
rect 8110 9568 8116 9580
rect 7883 9540 8116 9568
rect 7883 9537 7895 9540
rect 7837 9531 7895 9537
rect 5534 9460 5540 9512
rect 5592 9500 5598 9512
rect 6012 9500 6040 9531
rect 8110 9528 8116 9540
rect 8168 9528 8174 9580
rect 8573 9571 8631 9577
rect 8573 9568 8585 9571
rect 8220 9540 8585 9568
rect 5592 9472 6040 9500
rect 7285 9503 7343 9509
rect 5592 9460 5598 9472
rect 7285 9469 7297 9503
rect 7331 9500 7343 9503
rect 7374 9500 7380 9512
rect 7331 9472 7380 9500
rect 7331 9469 7343 9472
rect 7285 9463 7343 9469
rect 7374 9460 7380 9472
rect 7432 9460 7438 9512
rect 7561 9503 7619 9509
rect 7561 9469 7573 9503
rect 7607 9469 7619 9503
rect 7561 9463 7619 9469
rect 7929 9503 7987 9509
rect 7929 9469 7941 9503
rect 7975 9500 7987 9503
rect 8220 9500 8248 9540
rect 8573 9537 8585 9540
rect 8619 9568 8631 9571
rect 8662 9568 8668 9580
rect 8619 9540 8668 9568
rect 8619 9537 8631 9540
rect 8573 9531 8631 9537
rect 8662 9528 8668 9540
rect 8720 9528 8726 9580
rect 12802 9528 12808 9580
rect 12860 9528 12866 9580
rect 12897 9571 12955 9577
rect 12897 9537 12909 9571
rect 12943 9568 12955 9571
rect 13722 9568 13728 9580
rect 12943 9540 13728 9568
rect 12943 9537 12955 9540
rect 12897 9531 12955 9537
rect 13722 9528 13728 9540
rect 13780 9528 13786 9580
rect 15565 9571 15623 9577
rect 15565 9537 15577 9571
rect 15611 9537 15623 9571
rect 15565 9531 15623 9537
rect 15749 9571 15807 9577
rect 15749 9537 15761 9571
rect 15795 9568 15807 9571
rect 15930 9568 15936 9580
rect 15795 9540 15936 9568
rect 15795 9537 15807 9540
rect 15749 9531 15807 9537
rect 7975 9472 8248 9500
rect 7975 9469 7987 9472
rect 7929 9463 7987 9469
rect 7576 9432 7604 9463
rect 8294 9460 8300 9512
rect 8352 9460 8358 9512
rect 8478 9460 8484 9512
rect 8536 9460 8542 9512
rect 9122 9460 9128 9512
rect 9180 9460 9186 9512
rect 9401 9503 9459 9509
rect 9401 9500 9413 9503
rect 9232 9472 9413 9500
rect 8846 9432 8852 9444
rect 1636 9404 2774 9432
rect 2884 9404 3188 9432
rect 6104 9404 8852 9432
rect 1636 9392 1642 9404
rect 1486 9324 1492 9376
rect 1544 9324 1550 9376
rect 1670 9324 1676 9376
rect 1728 9364 1734 9376
rect 1765 9367 1823 9373
rect 1765 9364 1777 9367
rect 1728 9336 1777 9364
rect 1728 9324 1734 9336
rect 1765 9333 1777 9336
rect 1811 9333 1823 9367
rect 2746 9364 2774 9404
rect 6104 9364 6132 9404
rect 8846 9392 8852 9404
rect 8904 9392 8910 9444
rect 8941 9435 8999 9441
rect 8941 9401 8953 9435
rect 8987 9432 8999 9435
rect 9232 9432 9260 9472
rect 9401 9469 9413 9472
rect 9447 9469 9459 9503
rect 15580 9500 15608 9531
rect 15930 9528 15936 9540
rect 15988 9528 15994 9580
rect 16209 9571 16267 9577
rect 16209 9537 16221 9571
rect 16255 9568 16267 9571
rect 16298 9568 16304 9580
rect 16255 9540 16304 9568
rect 16255 9537 16267 9540
rect 16209 9531 16267 9537
rect 16298 9528 16304 9540
rect 16356 9528 16362 9580
rect 16485 9571 16543 9577
rect 16485 9537 16497 9571
rect 16531 9568 16543 9571
rect 16850 9568 16856 9580
rect 16531 9540 16856 9568
rect 16531 9537 16543 9540
rect 16485 9531 16543 9537
rect 16850 9528 16856 9540
rect 16908 9528 16914 9580
rect 16025 9503 16083 9509
rect 16025 9500 16037 9503
rect 15580 9472 16037 9500
rect 9401 9463 9459 9469
rect 16025 9469 16037 9472
rect 16071 9500 16083 9503
rect 16114 9500 16120 9512
rect 16071 9472 16120 9500
rect 16071 9469 16083 9472
rect 16025 9463 16083 9469
rect 16114 9460 16120 9472
rect 16172 9460 16178 9512
rect 8987 9404 9260 9432
rect 8987 9401 8999 9404
rect 8941 9395 8999 9401
rect 2746 9336 6132 9364
rect 6181 9367 6239 9373
rect 1765 9327 1823 9333
rect 6181 9333 6193 9367
rect 6227 9364 6239 9367
rect 6362 9364 6368 9376
rect 6227 9336 6368 9364
rect 6227 9333 6239 9336
rect 6181 9327 6239 9333
rect 6362 9324 6368 9336
rect 6420 9324 6426 9376
rect 6914 9324 6920 9376
rect 6972 9364 6978 9376
rect 7653 9367 7711 9373
rect 7653 9364 7665 9367
rect 6972 9336 7665 9364
rect 6972 9324 6978 9336
rect 7653 9333 7665 9336
rect 7699 9333 7711 9367
rect 7653 9327 7711 9333
rect 10686 9324 10692 9376
rect 10744 9364 10750 9376
rect 10873 9367 10931 9373
rect 10873 9364 10885 9367
rect 10744 9336 10885 9364
rect 10744 9324 10750 9336
rect 10873 9333 10885 9336
rect 10919 9333 10931 9367
rect 10873 9327 10931 9333
rect 1104 9274 17388 9296
rect 1104 9222 2985 9274
rect 3037 9222 3049 9274
rect 3101 9222 3113 9274
rect 3165 9222 3177 9274
rect 3229 9222 3241 9274
rect 3293 9222 7056 9274
rect 7108 9222 7120 9274
rect 7172 9222 7184 9274
rect 7236 9222 7248 9274
rect 7300 9222 7312 9274
rect 7364 9222 11127 9274
rect 11179 9222 11191 9274
rect 11243 9222 11255 9274
rect 11307 9222 11319 9274
rect 11371 9222 11383 9274
rect 11435 9222 15198 9274
rect 15250 9222 15262 9274
rect 15314 9222 15326 9274
rect 15378 9222 15390 9274
rect 15442 9222 15454 9274
rect 15506 9222 17388 9274
rect 1104 9200 17388 9222
rect 2682 9120 2688 9172
rect 2740 9160 2746 9172
rect 3145 9163 3203 9169
rect 3145 9160 3157 9163
rect 2740 9132 3157 9160
rect 2740 9120 2746 9132
rect 3145 9129 3157 9132
rect 3191 9129 3203 9163
rect 3145 9123 3203 9129
rect 1670 8984 1676 9036
rect 1728 8984 1734 9036
rect 1397 8959 1455 8965
rect 1397 8925 1409 8959
rect 1443 8925 1455 8959
rect 3160 8956 3188 9123
rect 3326 9120 3332 9172
rect 3384 9120 3390 9172
rect 7374 9160 7380 9172
rect 6656 9132 7380 9160
rect 6656 9033 6684 9132
rect 7374 9120 7380 9132
rect 7432 9120 7438 9172
rect 8294 9120 8300 9172
rect 8352 9160 8358 9172
rect 8573 9163 8631 9169
rect 8573 9160 8585 9163
rect 8352 9132 8585 9160
rect 8352 9120 8358 9132
rect 8573 9129 8585 9132
rect 8619 9129 8631 9163
rect 8573 9123 8631 9129
rect 15746 9120 15752 9172
rect 15804 9160 15810 9172
rect 15841 9163 15899 9169
rect 15841 9160 15853 9163
rect 15804 9132 15853 9160
rect 15804 9120 15810 9132
rect 15841 9129 15853 9132
rect 15887 9129 15899 9163
rect 15841 9123 15899 9129
rect 9122 9052 9128 9104
rect 9180 9092 9186 9104
rect 9217 9095 9275 9101
rect 9217 9092 9229 9095
rect 9180 9064 9229 9092
rect 9180 9052 9186 9064
rect 9217 9061 9229 9064
rect 9263 9061 9275 9095
rect 15856 9092 15884 9123
rect 15930 9120 15936 9172
rect 15988 9160 15994 9172
rect 15988 9132 16436 9160
rect 15988 9120 15994 9132
rect 16408 9092 16436 9132
rect 16761 9095 16819 9101
rect 16761 9092 16773 9095
rect 15856 9064 16252 9092
rect 9217 9055 9275 9061
rect 4065 9027 4123 9033
rect 4065 8993 4077 9027
rect 4111 9024 4123 9027
rect 5629 9027 5687 9033
rect 5629 9024 5641 9027
rect 4111 8996 5641 9024
rect 4111 8993 4123 8996
rect 4065 8987 4123 8993
rect 5629 8993 5641 8996
rect 5675 8993 5687 9027
rect 5629 8987 5687 8993
rect 5813 9027 5871 9033
rect 5813 8993 5825 9027
rect 5859 9024 5871 9027
rect 6641 9027 6699 9033
rect 5859 8996 6408 9024
rect 5859 8993 5871 8996
rect 5813 8987 5871 8993
rect 6380 8968 6408 8996
rect 6641 8993 6653 9027
rect 6687 8993 6699 9027
rect 6641 8987 6699 8993
rect 6914 8984 6920 9036
rect 6972 8984 6978 9036
rect 10594 8984 10600 9036
rect 10652 8984 10658 9036
rect 16114 8984 16120 9036
rect 16172 8984 16178 9036
rect 16224 9033 16252 9064
rect 16408 9064 16773 9092
rect 16209 9027 16267 9033
rect 16209 8993 16221 9027
rect 16255 8993 16267 9027
rect 16408 9024 16436 9064
rect 16761 9061 16773 9064
rect 16807 9061 16819 9095
rect 16761 9055 16819 9061
rect 16577 9027 16635 9033
rect 16577 9024 16589 9027
rect 16408 8996 16589 9024
rect 16209 8987 16267 8993
rect 16577 8993 16589 8996
rect 16623 8993 16635 9027
rect 16577 8987 16635 8993
rect 3237 8959 3295 8965
rect 3237 8956 3249 8959
rect 3160 8928 3249 8956
rect 1397 8919 1455 8925
rect 3237 8925 3249 8928
rect 3283 8925 3295 8959
rect 3237 8919 3295 8925
rect 1412 8888 1440 8919
rect 3418 8916 3424 8968
rect 3476 8916 3482 8968
rect 3510 8916 3516 8968
rect 3568 8916 3574 8968
rect 3789 8959 3847 8965
rect 3789 8925 3801 8959
rect 3835 8925 3847 8959
rect 3789 8919 3847 8925
rect 5905 8959 5963 8965
rect 5905 8925 5917 8959
rect 5951 8956 5963 8959
rect 6178 8956 6184 8968
rect 5951 8928 6184 8956
rect 5951 8925 5963 8928
rect 5905 8919 5963 8925
rect 3694 8888 3700 8900
rect 1412 8860 1624 8888
rect 2898 8860 3700 8888
rect 1596 8832 1624 8860
rect 3694 8848 3700 8860
rect 3752 8848 3758 8900
rect 1578 8780 1584 8832
rect 1636 8820 1642 8832
rect 3804 8820 3832 8919
rect 6178 8916 6184 8928
rect 6236 8916 6242 8968
rect 6362 8916 6368 8968
rect 6420 8916 6426 8968
rect 6546 8916 6552 8968
rect 6604 8916 6610 8968
rect 8754 8916 8760 8968
rect 8812 8916 8818 8968
rect 8846 8916 8852 8968
rect 8904 8956 8910 8968
rect 9401 8959 9459 8965
rect 9401 8956 9413 8959
rect 8904 8928 9413 8956
rect 8904 8916 8910 8928
rect 9401 8925 9413 8928
rect 9447 8925 9459 8959
rect 9401 8919 9459 8925
rect 5350 8888 5356 8900
rect 5290 8860 5356 8888
rect 5350 8848 5356 8860
rect 5408 8848 5414 8900
rect 6273 8891 6331 8897
rect 6273 8857 6285 8891
rect 6319 8888 6331 8891
rect 6564 8888 6592 8916
rect 6319 8860 6592 8888
rect 6319 8857 6331 8860
rect 6273 8851 6331 8857
rect 7374 8848 7380 8900
rect 7432 8848 7438 8900
rect 8481 8891 8539 8897
rect 8481 8857 8493 8891
rect 8527 8857 8539 8891
rect 8481 8851 8539 8857
rect 4706 8820 4712 8832
rect 1636 8792 4712 8820
rect 1636 8780 1642 8792
rect 4706 8780 4712 8792
rect 4764 8780 4770 8832
rect 5534 8780 5540 8832
rect 5592 8780 5598 8832
rect 6454 8780 6460 8832
rect 6512 8780 6518 8832
rect 8386 8780 8392 8832
rect 8444 8820 8450 8832
rect 8496 8820 8524 8851
rect 8662 8848 8668 8900
rect 8720 8848 8726 8900
rect 9416 8888 9444 8919
rect 10686 8916 10692 8968
rect 10744 8916 10750 8968
rect 13081 8959 13139 8965
rect 13081 8956 13093 8959
rect 12406 8928 13093 8956
rect 12406 8888 12434 8928
rect 13081 8925 13093 8928
rect 13127 8925 13139 8959
rect 13081 8919 13139 8925
rect 13357 8959 13415 8965
rect 13357 8925 13369 8959
rect 13403 8956 13415 8959
rect 14090 8956 14096 8968
rect 13403 8928 14096 8956
rect 13403 8925 13415 8928
rect 13357 8919 13415 8925
rect 14090 8916 14096 8928
rect 14148 8916 14154 8968
rect 15502 8928 16068 8956
rect 9416 8860 12434 8888
rect 13906 8848 13912 8900
rect 13964 8888 13970 8900
rect 14369 8891 14427 8897
rect 14369 8888 14381 8891
rect 13964 8860 14381 8888
rect 13964 8848 13970 8860
rect 14369 8857 14381 8860
rect 14415 8857 14427 8891
rect 15933 8891 15991 8897
rect 15933 8888 15945 8891
rect 14369 8851 14427 8857
rect 15672 8860 15945 8888
rect 8444 8792 8524 8820
rect 8444 8780 8450 8792
rect 11054 8780 11060 8832
rect 11112 8780 11118 8832
rect 15010 8780 15016 8832
rect 15068 8820 15074 8832
rect 15672 8820 15700 8860
rect 15933 8857 15945 8860
rect 15979 8857 15991 8891
rect 16040 8888 16068 8928
rect 16298 8916 16304 8968
rect 16356 8956 16362 8968
rect 16669 8959 16727 8965
rect 16669 8956 16681 8959
rect 16356 8928 16681 8956
rect 16356 8916 16362 8928
rect 16669 8925 16681 8928
rect 16715 8925 16727 8959
rect 16669 8919 16727 8925
rect 16850 8916 16856 8968
rect 16908 8916 16914 8968
rect 16942 8916 16948 8968
rect 17000 8916 17006 8968
rect 16390 8888 16396 8900
rect 16040 8860 16396 8888
rect 15933 8851 15991 8857
rect 16390 8848 16396 8860
rect 16448 8848 16454 8900
rect 15068 8792 15700 8820
rect 15068 8780 15074 8792
rect 1104 8730 17388 8752
rect 1104 8678 3645 8730
rect 3697 8678 3709 8730
rect 3761 8678 3773 8730
rect 3825 8678 3837 8730
rect 3889 8678 3901 8730
rect 3953 8678 7716 8730
rect 7768 8678 7780 8730
rect 7832 8678 7844 8730
rect 7896 8678 7908 8730
rect 7960 8678 7972 8730
rect 8024 8678 11787 8730
rect 11839 8678 11851 8730
rect 11903 8678 11915 8730
rect 11967 8678 11979 8730
rect 12031 8678 12043 8730
rect 12095 8678 15858 8730
rect 15910 8678 15922 8730
rect 15974 8678 15986 8730
rect 16038 8678 16050 8730
rect 16102 8678 16114 8730
rect 16166 8678 17388 8730
rect 1104 8656 17388 8678
rect 1857 8619 1915 8625
rect 1857 8585 1869 8619
rect 1903 8585 1915 8619
rect 1857 8579 1915 8585
rect 1872 8548 1900 8579
rect 2038 8576 2044 8628
rect 2096 8616 2102 8628
rect 2961 8619 3019 8625
rect 2961 8616 2973 8619
rect 2096 8588 2973 8616
rect 2096 8576 2102 8588
rect 2961 8585 2973 8588
rect 3007 8585 3019 8619
rect 5718 8616 5724 8628
rect 2961 8579 3019 8585
rect 3160 8588 5724 8616
rect 3160 8548 3188 8588
rect 5718 8576 5724 8588
rect 5776 8616 5782 8628
rect 5776 8588 6500 8616
rect 5776 8576 5782 8588
rect 1872 8520 3188 8548
rect 3970 8508 3976 8560
rect 4028 8508 4034 8560
rect 4433 8551 4491 8557
rect 4433 8517 4445 8551
rect 4479 8548 4491 8551
rect 4479 8520 5488 8548
rect 4479 8517 4491 8520
rect 4433 8511 4491 8517
rect 842 8440 848 8492
rect 900 8480 906 8492
rect 1397 8483 1455 8489
rect 1397 8480 1409 8483
rect 900 8452 1409 8480
rect 900 8440 906 8452
rect 1397 8449 1409 8452
rect 1443 8449 1455 8483
rect 1397 8443 1455 8449
rect 1670 8440 1676 8492
rect 1728 8440 1734 8492
rect 4706 8440 4712 8492
rect 4764 8440 4770 8492
rect 2746 8384 5396 8412
rect 1581 8347 1639 8353
rect 1581 8313 1593 8347
rect 1627 8344 1639 8347
rect 2746 8344 2774 8384
rect 1627 8316 2774 8344
rect 1627 8313 1639 8316
rect 1581 8307 1639 8313
rect 2406 8236 2412 8288
rect 2464 8276 2470 8288
rect 3418 8276 3424 8288
rect 2464 8248 3424 8276
rect 2464 8236 2470 8248
rect 3418 8236 3424 8248
rect 3476 8236 3482 8288
rect 3970 8236 3976 8288
rect 4028 8276 4034 8288
rect 5258 8276 5264 8288
rect 4028 8248 5264 8276
rect 4028 8236 4034 8248
rect 5258 8236 5264 8248
rect 5316 8236 5322 8288
rect 5368 8276 5396 8384
rect 5460 8353 5488 8520
rect 5534 8508 5540 8560
rect 5592 8548 5598 8560
rect 6365 8551 6423 8557
rect 6365 8548 6377 8551
rect 5592 8520 6377 8548
rect 5592 8508 5598 8520
rect 6365 8517 6377 8520
rect 6411 8517 6423 8551
rect 6365 8511 6423 8517
rect 5813 8483 5871 8489
rect 5813 8449 5825 8483
rect 5859 8480 5871 8483
rect 6178 8480 6184 8492
rect 5859 8452 6184 8480
rect 5859 8449 5871 8452
rect 5813 8443 5871 8449
rect 6178 8440 6184 8452
rect 6236 8440 6242 8492
rect 6472 8480 6500 8588
rect 6546 8576 6552 8628
rect 6604 8576 6610 8628
rect 7837 8619 7895 8625
rect 7837 8585 7849 8619
rect 7883 8616 7895 8619
rect 8110 8616 8116 8628
rect 7883 8588 8116 8616
rect 7883 8585 7895 8588
rect 7837 8579 7895 8585
rect 8110 8576 8116 8588
rect 8168 8576 8174 8628
rect 10594 8576 10600 8628
rect 10652 8576 10658 8628
rect 10686 8576 10692 8628
rect 10744 8576 10750 8628
rect 13906 8576 13912 8628
rect 13964 8576 13970 8628
rect 16298 8576 16304 8628
rect 16356 8616 16362 8628
rect 16485 8619 16543 8625
rect 16485 8616 16497 8619
rect 16356 8588 16497 8616
rect 16356 8576 16362 8588
rect 16485 8585 16497 8588
rect 16531 8585 16543 8619
rect 16485 8579 16543 8585
rect 16850 8576 16856 8628
rect 16908 8576 16914 8628
rect 8386 8548 8392 8560
rect 8036 8520 8392 8548
rect 6549 8483 6607 8489
rect 6549 8480 6561 8483
rect 6472 8452 6561 8480
rect 6549 8449 6561 8452
rect 6595 8449 6607 8483
rect 6549 8443 6607 8449
rect 6641 8483 6699 8489
rect 6641 8449 6653 8483
rect 6687 8480 6699 8483
rect 6730 8480 6736 8492
rect 6687 8452 6736 8480
rect 6687 8449 6699 8452
rect 6641 8443 6699 8449
rect 6730 8440 6736 8452
rect 6788 8440 6794 8492
rect 8036 8489 8064 8520
rect 8386 8508 8392 8520
rect 8444 8508 8450 8560
rect 10704 8548 10732 8576
rect 10060 8520 10732 8548
rect 8021 8483 8079 8489
rect 8021 8449 8033 8483
rect 8067 8449 8079 8483
rect 8021 8443 8079 8449
rect 8205 8483 8263 8489
rect 8205 8449 8217 8483
rect 8251 8449 8263 8483
rect 8205 8443 8263 8449
rect 8297 8483 8355 8489
rect 8297 8449 8309 8483
rect 8343 8480 8355 8483
rect 8662 8480 8668 8492
rect 8343 8452 8668 8480
rect 8343 8449 8355 8452
rect 8297 8443 8355 8449
rect 5905 8415 5963 8421
rect 5905 8381 5917 8415
rect 5951 8412 5963 8415
rect 6454 8412 6460 8424
rect 5951 8384 6460 8412
rect 5951 8381 5963 8384
rect 5905 8375 5963 8381
rect 6454 8372 6460 8384
rect 6512 8372 6518 8424
rect 6914 8372 6920 8424
rect 6972 8412 6978 8424
rect 7558 8412 7564 8424
rect 6972 8384 7564 8412
rect 6972 8372 6978 8384
rect 7558 8372 7564 8384
rect 7616 8412 7622 8424
rect 8220 8412 8248 8443
rect 7616 8384 8248 8412
rect 7616 8372 7622 8384
rect 5445 8347 5503 8353
rect 5445 8313 5457 8347
rect 5491 8313 5503 8347
rect 8312 8344 8340 8443
rect 8662 8440 8668 8452
rect 8720 8440 8726 8492
rect 10060 8489 10088 8520
rect 11054 8508 11060 8560
rect 11112 8548 11118 8560
rect 11793 8551 11851 8557
rect 11793 8548 11805 8551
rect 11112 8520 11805 8548
rect 11112 8508 11118 8520
rect 11793 8517 11805 8520
rect 11839 8517 11851 8551
rect 11793 8511 11851 8517
rect 12434 8508 12440 8560
rect 12492 8508 12498 8560
rect 15010 8508 15016 8560
rect 15068 8508 15074 8560
rect 16390 8548 16396 8560
rect 16238 8520 16396 8548
rect 16390 8508 16396 8520
rect 16448 8508 16454 8560
rect 10045 8483 10103 8489
rect 10045 8449 10057 8483
rect 10091 8449 10103 8483
rect 10045 8443 10103 8449
rect 10505 8483 10563 8489
rect 10505 8449 10517 8483
rect 10551 8449 10563 8483
rect 10505 8443 10563 8449
rect 10689 8483 10747 8489
rect 10689 8449 10701 8483
rect 10735 8449 10747 8483
rect 13541 8483 13599 8489
rect 13541 8480 13553 8483
rect 10689 8443 10747 8449
rect 13280 8452 13553 8480
rect 9953 8415 10011 8421
rect 9953 8381 9965 8415
rect 9999 8381 10011 8415
rect 9953 8375 10011 8381
rect 5445 8307 5503 8313
rect 5552 8316 8340 8344
rect 9968 8344 9996 8375
rect 10410 8372 10416 8424
rect 10468 8412 10474 8424
rect 10520 8412 10548 8443
rect 10468 8384 10548 8412
rect 10468 8372 10474 8384
rect 10704 8344 10732 8443
rect 11514 8372 11520 8424
rect 11572 8372 11578 8424
rect 13280 8421 13308 8452
rect 13541 8449 13553 8452
rect 13587 8480 13599 8483
rect 13630 8480 13636 8492
rect 13587 8452 13636 8480
rect 13587 8449 13599 8452
rect 13541 8443 13599 8449
rect 13630 8440 13636 8452
rect 13688 8440 13694 8492
rect 14090 8440 14096 8492
rect 14148 8480 14154 8492
rect 14550 8480 14556 8492
rect 14148 8452 14556 8480
rect 14148 8440 14154 8452
rect 14550 8440 14556 8452
rect 14608 8480 14614 8492
rect 14737 8483 14795 8489
rect 14737 8480 14749 8483
rect 14608 8452 14749 8480
rect 14608 8440 14614 8452
rect 14737 8449 14749 8452
rect 14783 8449 14795 8483
rect 14737 8443 14795 8449
rect 17034 8440 17040 8492
rect 17092 8440 17098 8492
rect 13265 8415 13323 8421
rect 13265 8381 13277 8415
rect 13311 8381 13323 8415
rect 13265 8375 13323 8381
rect 13446 8372 13452 8424
rect 13504 8372 13510 8424
rect 10778 8344 10784 8356
rect 9968 8316 10784 8344
rect 5552 8276 5580 8316
rect 10778 8304 10784 8316
rect 10836 8304 10842 8356
rect 5368 8248 5580 8276
rect 9766 8236 9772 8288
rect 9824 8236 9830 8288
rect 1104 8186 17388 8208
rect 1104 8134 2985 8186
rect 3037 8134 3049 8186
rect 3101 8134 3113 8186
rect 3165 8134 3177 8186
rect 3229 8134 3241 8186
rect 3293 8134 7056 8186
rect 7108 8134 7120 8186
rect 7172 8134 7184 8186
rect 7236 8134 7248 8186
rect 7300 8134 7312 8186
rect 7364 8134 11127 8186
rect 11179 8134 11191 8186
rect 11243 8134 11255 8186
rect 11307 8134 11319 8186
rect 11371 8134 11383 8186
rect 11435 8134 15198 8186
rect 15250 8134 15262 8186
rect 15314 8134 15326 8186
rect 15378 8134 15390 8186
rect 15442 8134 15454 8186
rect 15506 8134 17388 8186
rect 1104 8112 17388 8134
rect 1581 8075 1639 8081
rect 1581 8041 1593 8075
rect 1627 8072 1639 8075
rect 2222 8072 2228 8084
rect 1627 8044 2228 8072
rect 1627 8041 1639 8044
rect 1581 8035 1639 8041
rect 2222 8032 2228 8044
rect 2280 8072 2286 8084
rect 3329 8075 3387 8081
rect 3329 8072 3341 8075
rect 2280 8044 3341 8072
rect 2280 8032 2286 8044
rect 3329 8041 3341 8044
rect 3375 8041 3387 8075
rect 3329 8035 3387 8041
rect 10778 8032 10784 8084
rect 10836 8032 10842 8084
rect 13265 8075 13323 8081
rect 13265 8041 13277 8075
rect 13311 8072 13323 8075
rect 13446 8072 13452 8084
rect 13311 8044 13452 8072
rect 13311 8041 13323 8044
rect 13265 8035 13323 8041
rect 13446 8032 13452 8044
rect 13504 8032 13510 8084
rect 8202 8004 8208 8016
rect 7668 7976 8208 8004
rect 842 7828 848 7880
rect 900 7868 906 7880
rect 7668 7877 7696 7976
rect 8202 7964 8208 7976
rect 8260 8004 8266 8016
rect 8662 8004 8668 8016
rect 8260 7976 8668 8004
rect 8260 7964 8266 7976
rect 8662 7964 8668 7976
rect 8720 7964 8726 8016
rect 8294 7936 8300 7948
rect 7760 7908 8300 7936
rect 7760 7877 7788 7908
rect 8294 7896 8300 7908
rect 8352 7896 8358 7948
rect 9217 7939 9275 7945
rect 9217 7905 9229 7939
rect 9263 7936 9275 7939
rect 9766 7936 9772 7948
rect 9263 7908 9772 7936
rect 9263 7905 9275 7908
rect 9217 7899 9275 7905
rect 9766 7896 9772 7908
rect 9824 7896 9830 7948
rect 1397 7871 1455 7877
rect 1397 7868 1409 7871
rect 900 7840 1409 7868
rect 900 7828 906 7840
rect 1397 7837 1409 7840
rect 1443 7837 1455 7871
rect 1397 7831 1455 7837
rect 7653 7871 7711 7877
rect 7653 7837 7665 7871
rect 7699 7837 7711 7871
rect 7653 7831 7711 7837
rect 7745 7871 7803 7877
rect 7745 7837 7757 7871
rect 7791 7837 7803 7871
rect 8021 7871 8079 7877
rect 8021 7868 8033 7871
rect 7745 7831 7803 7837
rect 7852 7840 8033 7868
rect 3513 7803 3571 7809
rect 3513 7769 3525 7803
rect 3559 7800 3571 7803
rect 6914 7800 6920 7812
rect 3559 7772 6920 7800
rect 3559 7769 3571 7772
rect 3513 7763 3571 7769
rect 6914 7760 6920 7772
rect 6972 7760 6978 7812
rect 3142 7692 3148 7744
rect 3200 7692 3206 7744
rect 3313 7735 3371 7741
rect 3313 7701 3325 7735
rect 3359 7732 3371 7735
rect 3418 7732 3424 7744
rect 3359 7704 3424 7732
rect 3359 7701 3371 7704
rect 3313 7695 3371 7701
rect 3418 7692 3424 7704
rect 3476 7692 3482 7744
rect 7558 7692 7564 7744
rect 7616 7732 7622 7744
rect 7653 7735 7711 7741
rect 7653 7732 7665 7735
rect 7616 7704 7665 7732
rect 7616 7692 7622 7704
rect 7653 7701 7665 7704
rect 7699 7732 7711 7735
rect 7852 7732 7880 7840
rect 8021 7837 8033 7840
rect 8067 7837 8079 7871
rect 8021 7831 8079 7837
rect 8202 7828 8208 7880
rect 8260 7828 8266 7880
rect 8941 7871 8999 7877
rect 8941 7837 8953 7871
rect 8987 7837 8999 7871
rect 10965 7871 11023 7877
rect 10965 7868 10977 7871
rect 8941 7831 8999 7837
rect 10704 7840 10977 7868
rect 7929 7803 7987 7809
rect 7929 7769 7941 7803
rect 7975 7800 7987 7803
rect 8110 7800 8116 7812
rect 7975 7772 8116 7800
rect 7975 7769 7987 7772
rect 7929 7763 7987 7769
rect 8110 7760 8116 7772
rect 8168 7760 8174 7812
rect 8956 7800 8984 7831
rect 9122 7800 9128 7812
rect 8956 7772 9128 7800
rect 9122 7760 9128 7772
rect 9180 7760 9186 7812
rect 9950 7760 9956 7812
rect 10008 7760 10014 7812
rect 10704 7744 10732 7840
rect 10965 7837 10977 7840
rect 11011 7837 11023 7871
rect 10965 7831 11023 7837
rect 11241 7871 11299 7877
rect 11241 7837 11253 7871
rect 11287 7837 11299 7871
rect 11241 7831 11299 7837
rect 13173 7871 13231 7877
rect 13173 7837 13185 7871
rect 13219 7837 13231 7871
rect 13173 7831 13231 7837
rect 13357 7871 13415 7877
rect 13357 7837 13369 7871
rect 13403 7868 13415 7871
rect 13538 7868 13544 7880
rect 13403 7840 13544 7868
rect 13403 7837 13415 7840
rect 13357 7831 13415 7837
rect 10870 7760 10876 7812
rect 10928 7800 10934 7812
rect 11256 7800 11284 7831
rect 10928 7772 11284 7800
rect 13188 7800 13216 7831
rect 13538 7828 13544 7840
rect 13596 7828 13602 7880
rect 17034 7828 17040 7880
rect 17092 7828 17098 7880
rect 13998 7800 14004 7812
rect 13188 7772 14004 7800
rect 10928 7760 10934 7772
rect 13998 7760 14004 7772
rect 14056 7760 14062 7812
rect 7699 7704 7880 7732
rect 8205 7735 8263 7741
rect 7699 7701 7711 7704
rect 7653 7695 7711 7701
rect 8205 7701 8217 7735
rect 8251 7732 8263 7735
rect 8478 7732 8484 7744
rect 8251 7704 8484 7732
rect 8251 7701 8263 7704
rect 8205 7695 8263 7701
rect 8478 7692 8484 7704
rect 8536 7692 8542 7744
rect 10686 7692 10692 7744
rect 10744 7692 10750 7744
rect 11149 7735 11207 7741
rect 11149 7701 11161 7735
rect 11195 7732 11207 7735
rect 12710 7732 12716 7744
rect 11195 7704 12716 7732
rect 11195 7701 11207 7704
rect 11149 7695 11207 7701
rect 12710 7692 12716 7704
rect 12768 7692 12774 7744
rect 14274 7692 14280 7744
rect 14332 7732 14338 7744
rect 16853 7735 16911 7741
rect 16853 7732 16865 7735
rect 14332 7704 16865 7732
rect 14332 7692 14338 7704
rect 16853 7701 16865 7704
rect 16899 7701 16911 7735
rect 16853 7695 16911 7701
rect 1104 7642 17388 7664
rect 1104 7590 3645 7642
rect 3697 7590 3709 7642
rect 3761 7590 3773 7642
rect 3825 7590 3837 7642
rect 3889 7590 3901 7642
rect 3953 7590 7716 7642
rect 7768 7590 7780 7642
rect 7832 7590 7844 7642
rect 7896 7590 7908 7642
rect 7960 7590 7972 7642
rect 8024 7590 11787 7642
rect 11839 7590 11851 7642
rect 11903 7590 11915 7642
rect 11967 7590 11979 7642
rect 12031 7590 12043 7642
rect 12095 7590 15858 7642
rect 15910 7590 15922 7642
rect 15974 7590 15986 7642
rect 16038 7590 16050 7642
rect 16102 7590 16114 7642
rect 16166 7590 17388 7642
rect 1104 7568 17388 7590
rect 6178 7488 6184 7540
rect 6236 7488 6242 7540
rect 7374 7488 7380 7540
rect 7432 7528 7438 7540
rect 7650 7528 7656 7540
rect 7432 7500 7656 7528
rect 7432 7488 7438 7500
rect 7650 7488 7656 7500
rect 7708 7488 7714 7540
rect 8110 7488 8116 7540
rect 8168 7488 8174 7540
rect 10045 7531 10103 7537
rect 10045 7497 10057 7531
rect 10091 7528 10103 7531
rect 10410 7528 10416 7540
rect 10091 7500 10416 7528
rect 10091 7497 10103 7500
rect 10045 7491 10103 7497
rect 10410 7488 10416 7500
rect 10468 7488 10474 7540
rect 13265 7531 13323 7537
rect 13265 7497 13277 7531
rect 13311 7497 13323 7531
rect 13265 7491 13323 7497
rect 3602 7420 3608 7472
rect 3660 7460 3666 7472
rect 3970 7460 3976 7472
rect 3660 7432 3976 7460
rect 3660 7420 3666 7432
rect 3970 7420 3976 7432
rect 4028 7420 4034 7472
rect 4706 7460 4712 7472
rect 4448 7432 4712 7460
rect 2222 7352 2228 7404
rect 2280 7352 2286 7404
rect 2317 7395 2375 7401
rect 2317 7361 2329 7395
rect 2363 7392 2375 7395
rect 2406 7392 2412 7404
rect 2363 7364 2412 7392
rect 2363 7361 2375 7364
rect 2317 7355 2375 7361
rect 2406 7352 2412 7364
rect 2464 7352 2470 7404
rect 4448 7401 4476 7432
rect 4706 7420 4712 7432
rect 4764 7420 4770 7472
rect 5258 7420 5264 7472
rect 5316 7420 5322 7472
rect 6641 7463 6699 7469
rect 6641 7429 6653 7463
rect 6687 7460 6699 7463
rect 6914 7460 6920 7472
rect 6687 7432 6920 7460
rect 6687 7429 6699 7432
rect 6641 7423 6699 7429
rect 6914 7420 6920 7432
rect 6972 7420 6978 7472
rect 7282 7420 7288 7472
rect 7340 7420 7346 7472
rect 10137 7463 10195 7469
rect 10137 7429 10149 7463
rect 10183 7460 10195 7463
rect 10686 7460 10692 7472
rect 10183 7432 10692 7460
rect 10183 7429 10195 7432
rect 10137 7423 10195 7429
rect 10686 7420 10692 7432
rect 10744 7420 10750 7472
rect 12434 7420 12440 7472
rect 12492 7420 12498 7472
rect 13280 7460 13308 7491
rect 13998 7488 14004 7540
rect 14056 7528 14062 7540
rect 14185 7531 14243 7537
rect 14185 7528 14197 7531
rect 14056 7500 14197 7528
rect 14056 7488 14062 7500
rect 14185 7497 14197 7500
rect 14231 7497 14243 7531
rect 14185 7491 14243 7497
rect 13446 7460 13452 7472
rect 13280 7432 13452 7460
rect 13446 7420 13452 7432
rect 13504 7460 13510 7472
rect 14093 7463 14151 7469
rect 14093 7460 14105 7463
rect 13504 7432 14105 7460
rect 13504 7420 13510 7432
rect 14093 7429 14105 7432
rect 14139 7429 14151 7463
rect 14093 7423 14151 7429
rect 14274 7420 14280 7472
rect 14332 7420 14338 7472
rect 16390 7460 16396 7472
rect 16054 7432 16396 7460
rect 16390 7420 16396 7432
rect 16448 7420 16454 7472
rect 2501 7395 2559 7401
rect 2501 7361 2513 7395
rect 2547 7392 2559 7395
rect 4341 7395 4399 7401
rect 2547 7364 2774 7392
rect 2547 7361 2559 7364
rect 2501 7355 2559 7361
rect 2746 7324 2774 7364
rect 4341 7361 4353 7395
rect 4387 7392 4399 7395
rect 4433 7395 4491 7401
rect 4433 7392 4445 7395
rect 4387 7364 4445 7392
rect 4387 7361 4399 7364
rect 4341 7355 4399 7361
rect 4433 7361 4445 7364
rect 4479 7361 4491 7395
rect 4433 7355 4491 7361
rect 8018 7352 8024 7404
rect 8076 7392 8082 7404
rect 8573 7395 8631 7401
rect 8573 7392 8585 7395
rect 8076 7364 8585 7392
rect 8076 7352 8082 7364
rect 8573 7361 8585 7364
rect 8619 7361 8631 7395
rect 8573 7355 8631 7361
rect 8662 7352 8668 7404
rect 8720 7392 8726 7404
rect 9861 7395 9919 7401
rect 9861 7392 9873 7395
rect 8720 7364 9873 7392
rect 8720 7352 8726 7364
rect 9861 7361 9873 7364
rect 9907 7361 9919 7395
rect 9861 7355 9919 7361
rect 9953 7395 10011 7401
rect 9953 7361 9965 7395
rect 9999 7392 10011 7395
rect 10318 7392 10324 7404
rect 9999 7364 10324 7392
rect 9999 7361 10011 7364
rect 9953 7355 10011 7361
rect 10318 7352 10324 7364
rect 10376 7392 10382 7404
rect 10870 7392 10876 7404
rect 10376 7364 10876 7392
rect 10376 7352 10382 7364
rect 10870 7352 10876 7364
rect 10928 7352 10934 7404
rect 13630 7352 13636 7404
rect 13688 7352 13694 7404
rect 13814 7352 13820 7404
rect 13872 7392 13878 7404
rect 14369 7395 14427 7401
rect 14369 7392 14381 7395
rect 13872 7364 14381 7392
rect 13872 7352 13878 7364
rect 14369 7361 14381 7364
rect 14415 7361 14427 7395
rect 14369 7355 14427 7361
rect 14550 7352 14556 7404
rect 14608 7352 14614 7404
rect 17034 7352 17040 7404
rect 17092 7352 17098 7404
rect 3418 7324 3424 7336
rect 2746 7296 3424 7324
rect 3418 7284 3424 7296
rect 3476 7284 3482 7336
rect 4062 7284 4068 7336
rect 4120 7284 4126 7336
rect 4709 7327 4767 7333
rect 4709 7293 4721 7327
rect 4755 7324 4767 7327
rect 6365 7327 6423 7333
rect 4755 7296 6316 7324
rect 4755 7293 4767 7296
rect 4709 7287 4767 7293
rect 2501 7259 2559 7265
rect 2501 7225 2513 7259
rect 2547 7256 2559 7259
rect 2547 7228 3096 7256
rect 2547 7225 2559 7228
rect 2501 7219 2559 7225
rect 2593 7191 2651 7197
rect 2593 7157 2605 7191
rect 2639 7188 2651 7191
rect 2866 7188 2872 7200
rect 2639 7160 2872 7188
rect 2639 7157 2651 7160
rect 2593 7151 2651 7157
rect 2866 7148 2872 7160
rect 2924 7148 2930 7200
rect 3068 7188 3096 7228
rect 3970 7188 3976 7200
rect 3068 7160 3976 7188
rect 3970 7148 3976 7160
rect 4028 7148 4034 7200
rect 6288 7188 6316 7296
rect 6365 7293 6377 7327
rect 6411 7324 6423 7327
rect 7374 7324 7380 7336
rect 6411 7296 7380 7324
rect 6411 7293 6423 7296
rect 6365 7287 6423 7293
rect 7374 7284 7380 7296
rect 7432 7284 7438 7336
rect 8478 7284 8484 7336
rect 8536 7284 8542 7336
rect 9122 7284 9128 7336
rect 9180 7324 9186 7336
rect 11514 7324 11520 7336
rect 9180 7296 11520 7324
rect 9180 7284 9186 7296
rect 11514 7284 11520 7296
rect 11572 7284 11578 7336
rect 11793 7327 11851 7333
rect 11793 7293 11805 7327
rect 11839 7324 11851 7327
rect 13357 7327 13415 7333
rect 13357 7324 13369 7327
rect 11839 7296 13369 7324
rect 11839 7293 11851 7296
rect 11793 7287 11851 7293
rect 13357 7293 13369 7296
rect 13403 7293 13415 7327
rect 13357 7287 13415 7293
rect 13538 7284 13544 7336
rect 13596 7284 13602 7336
rect 14829 7327 14887 7333
rect 14829 7293 14841 7327
rect 14875 7324 14887 7327
rect 15562 7324 15568 7336
rect 14875 7296 15568 7324
rect 14875 7293 14887 7296
rect 14829 7287 14887 7293
rect 15562 7284 15568 7296
rect 15620 7284 15626 7336
rect 8205 7259 8263 7265
rect 8205 7225 8217 7259
rect 8251 7225 8263 7259
rect 8205 7219 8263 7225
rect 8220 7188 8248 7219
rect 6288 7160 8248 7188
rect 16298 7148 16304 7200
rect 16356 7148 16362 7200
rect 16666 7148 16672 7200
rect 16724 7188 16730 7200
rect 16853 7191 16911 7197
rect 16853 7188 16865 7191
rect 16724 7160 16865 7188
rect 16724 7148 16730 7160
rect 16853 7157 16865 7160
rect 16899 7157 16911 7191
rect 16853 7151 16911 7157
rect 1104 7098 17388 7120
rect 1104 7046 2985 7098
rect 3037 7046 3049 7098
rect 3101 7046 3113 7098
rect 3165 7046 3177 7098
rect 3229 7046 3241 7098
rect 3293 7046 7056 7098
rect 7108 7046 7120 7098
rect 7172 7046 7184 7098
rect 7236 7046 7248 7098
rect 7300 7046 7312 7098
rect 7364 7046 11127 7098
rect 11179 7046 11191 7098
rect 11243 7046 11255 7098
rect 11307 7046 11319 7098
rect 11371 7046 11383 7098
rect 11435 7046 15198 7098
rect 15250 7046 15262 7098
rect 15314 7046 15326 7098
rect 15378 7046 15390 7098
rect 15442 7046 15454 7098
rect 15506 7046 17388 7098
rect 1104 7024 17388 7046
rect 1660 6987 1718 6993
rect 1660 6953 1672 6987
rect 1706 6984 1718 6987
rect 3421 6987 3479 6993
rect 3421 6984 3433 6987
rect 1706 6956 3433 6984
rect 1706 6953 1718 6956
rect 1660 6947 1718 6953
rect 3421 6953 3433 6956
rect 3467 6953 3479 6987
rect 3421 6947 3479 6953
rect 3973 6987 4031 6993
rect 3973 6953 3985 6987
rect 4019 6984 4031 6987
rect 4062 6984 4068 6996
rect 4019 6956 4068 6984
rect 4019 6953 4031 6956
rect 3973 6947 4031 6953
rect 1397 6783 1455 6789
rect 1397 6749 1409 6783
rect 1443 6749 1455 6783
rect 1397 6743 1455 6749
rect 3237 6783 3295 6789
rect 3237 6749 3249 6783
rect 3283 6780 3295 6783
rect 3326 6780 3332 6792
rect 3283 6752 3332 6780
rect 3283 6749 3295 6752
rect 3237 6743 3295 6749
rect 1412 6712 1440 6743
rect 3326 6740 3332 6752
rect 3384 6740 3390 6792
rect 3436 6780 3464 6947
rect 4062 6944 4068 6956
rect 4120 6944 4126 6996
rect 7837 6987 7895 6993
rect 7837 6953 7849 6987
rect 7883 6984 7895 6987
rect 8202 6984 8208 6996
rect 7883 6956 8208 6984
rect 7883 6953 7895 6956
rect 7837 6947 7895 6953
rect 7852 6916 7880 6947
rect 8202 6944 8208 6956
rect 8260 6944 8266 6996
rect 13357 6987 13415 6993
rect 13357 6953 13369 6987
rect 13403 6984 13415 6987
rect 13538 6984 13544 6996
rect 13403 6956 13544 6984
rect 13403 6953 13415 6956
rect 13357 6947 13415 6953
rect 13538 6944 13544 6956
rect 13596 6944 13602 6996
rect 7300 6888 7880 6916
rect 16577 6919 16635 6925
rect 6914 6808 6920 6860
rect 6972 6848 6978 6860
rect 7300 6857 7328 6888
rect 16577 6885 16589 6919
rect 16623 6885 16635 6919
rect 16577 6879 16635 6885
rect 7101 6851 7159 6857
rect 7101 6848 7113 6851
rect 6972 6820 7113 6848
rect 6972 6808 6978 6820
rect 7101 6817 7113 6820
rect 7147 6817 7159 6851
rect 7101 6811 7159 6817
rect 7285 6851 7343 6857
rect 7285 6817 7297 6851
rect 7331 6817 7343 6851
rect 7285 6811 7343 6817
rect 7558 6808 7564 6860
rect 7616 6848 7622 6860
rect 7745 6851 7803 6857
rect 7745 6848 7757 6851
rect 7616 6820 7757 6848
rect 7616 6808 7622 6820
rect 7745 6817 7757 6820
rect 7791 6817 7803 6851
rect 7745 6811 7803 6817
rect 15197 6851 15255 6857
rect 15197 6817 15209 6851
rect 15243 6848 15255 6851
rect 15562 6848 15568 6860
rect 15243 6820 15568 6848
rect 15243 6817 15255 6820
rect 15197 6811 15255 6817
rect 15562 6808 15568 6820
rect 15620 6808 15626 6860
rect 15841 6851 15899 6857
rect 15841 6817 15853 6851
rect 15887 6848 15899 6851
rect 16206 6848 16212 6860
rect 15887 6820 16212 6848
rect 15887 6817 15899 6820
rect 15841 6811 15899 6817
rect 16206 6808 16212 6820
rect 16264 6848 16270 6860
rect 16592 6848 16620 6879
rect 16264 6820 16620 6848
rect 16264 6808 16270 6820
rect 3789 6783 3847 6789
rect 3789 6780 3801 6783
rect 3436 6752 3801 6780
rect 3789 6749 3801 6752
rect 3835 6749 3847 6783
rect 3789 6743 3847 6749
rect 3970 6740 3976 6792
rect 4028 6740 4034 6792
rect 4062 6740 4068 6792
rect 4120 6780 4126 6792
rect 5445 6783 5503 6789
rect 5445 6780 5457 6783
rect 4120 6752 5457 6780
rect 4120 6740 4126 6752
rect 5445 6749 5457 6752
rect 5491 6749 5503 6783
rect 5445 6743 5503 6749
rect 7377 6783 7435 6789
rect 7377 6749 7389 6783
rect 7423 6749 7435 6783
rect 7377 6743 7435 6749
rect 8021 6783 8079 6789
rect 8021 6749 8033 6783
rect 8067 6780 8079 6783
rect 8110 6780 8116 6792
rect 8067 6752 8116 6780
rect 8067 6749 8079 6752
rect 8021 6743 8079 6749
rect 1578 6712 1584 6724
rect 1412 6684 1584 6712
rect 1578 6672 1584 6684
rect 1636 6672 1642 6724
rect 3602 6712 3608 6724
rect 2898 6684 3608 6712
rect 3602 6672 3608 6684
rect 3660 6672 3666 6724
rect 4985 6715 5043 6721
rect 4985 6681 4997 6715
rect 5031 6712 5043 6715
rect 6181 6715 6239 6721
rect 6181 6712 6193 6715
rect 5031 6684 6193 6712
rect 5031 6681 5043 6684
rect 4985 6675 5043 6681
rect 3145 6647 3203 6653
rect 3145 6613 3157 6647
rect 3191 6644 3203 6647
rect 3418 6644 3424 6656
rect 3191 6616 3424 6644
rect 3191 6613 3203 6616
rect 3145 6607 3203 6613
rect 3418 6604 3424 6616
rect 3476 6604 3482 6656
rect 5074 6604 5080 6656
rect 5132 6604 5138 6656
rect 5644 6653 5672 6684
rect 6181 6681 6193 6684
rect 6227 6712 6239 6715
rect 6914 6712 6920 6724
rect 6227 6684 6920 6712
rect 6227 6681 6239 6684
rect 6181 6675 6239 6681
rect 6914 6672 6920 6684
rect 6972 6672 6978 6724
rect 5629 6647 5687 6653
rect 5629 6613 5641 6647
rect 5675 6613 5687 6647
rect 5629 6607 5687 6613
rect 5810 6604 5816 6656
rect 5868 6644 5874 6656
rect 6454 6644 6460 6656
rect 5868 6616 6460 6644
rect 5868 6604 5874 6616
rect 6454 6604 6460 6616
rect 6512 6604 6518 6656
rect 7392 6644 7420 6743
rect 8110 6740 8116 6752
rect 8168 6740 8174 6792
rect 8294 6740 8300 6792
rect 8352 6740 8358 6792
rect 13446 6740 13452 6792
rect 13504 6780 13510 6792
rect 13541 6783 13599 6789
rect 13541 6780 13553 6783
rect 13504 6752 13553 6780
rect 13504 6740 13510 6752
rect 13541 6749 13553 6752
rect 13587 6749 13599 6783
rect 13541 6743 13599 6749
rect 13722 6740 13728 6792
rect 13780 6740 13786 6792
rect 13817 6783 13875 6789
rect 13817 6749 13829 6783
rect 13863 6780 13875 6783
rect 14274 6780 14280 6792
rect 13863 6752 14280 6780
rect 13863 6749 13875 6752
rect 13817 6743 13875 6749
rect 14274 6740 14280 6752
rect 14332 6740 14338 6792
rect 15381 6783 15439 6789
rect 15381 6749 15393 6783
rect 15427 6749 15439 6783
rect 15381 6743 15439 6749
rect 15473 6783 15531 6789
rect 15473 6749 15485 6783
rect 15519 6780 15531 6783
rect 15654 6780 15660 6792
rect 15519 6752 15660 6780
rect 15519 6749 15531 6752
rect 15473 6743 15531 6749
rect 10962 6672 10968 6724
rect 11020 6712 11026 6724
rect 12802 6712 12808 6724
rect 11020 6684 12808 6712
rect 11020 6672 11026 6684
rect 12802 6672 12808 6684
rect 12860 6712 12866 6724
rect 13740 6712 13768 6740
rect 12860 6684 13768 6712
rect 15396 6712 15424 6743
rect 15654 6740 15660 6752
rect 15712 6740 15718 6792
rect 16117 6783 16175 6789
rect 16117 6749 16129 6783
rect 16163 6780 16175 6783
rect 16298 6780 16304 6792
rect 16163 6752 16304 6780
rect 16163 6749 16175 6752
rect 16117 6743 16175 6749
rect 16298 6740 16304 6752
rect 16356 6740 16362 6792
rect 16393 6783 16451 6789
rect 16393 6749 16405 6783
rect 16439 6780 16451 6783
rect 16666 6780 16672 6792
rect 16439 6752 16672 6780
rect 16439 6749 16451 6752
rect 16393 6743 16451 6749
rect 16666 6740 16672 6752
rect 16724 6740 16730 6792
rect 16761 6783 16819 6789
rect 16761 6749 16773 6783
rect 16807 6780 16819 6783
rect 16850 6780 16856 6792
rect 16807 6752 16856 6780
rect 16807 6749 16819 6752
rect 16761 6743 16819 6749
rect 16850 6740 16856 6752
rect 16908 6740 16914 6792
rect 15746 6712 15752 6724
rect 15396 6684 15752 6712
rect 12860 6672 12866 6684
rect 15746 6672 15752 6684
rect 15804 6712 15810 6724
rect 15933 6715 15991 6721
rect 15933 6712 15945 6715
rect 15804 6684 15945 6712
rect 15804 6672 15810 6684
rect 15933 6681 15945 6684
rect 15979 6681 15991 6715
rect 16316 6712 16344 6740
rect 16485 6715 16543 6721
rect 16485 6712 16497 6715
rect 16316 6684 16497 6712
rect 15933 6675 15991 6681
rect 16485 6681 16497 6684
rect 16531 6681 16543 6715
rect 16485 6675 16543 6681
rect 8110 6644 8116 6656
rect 7392 6616 8116 6644
rect 8110 6604 8116 6616
rect 8168 6604 8174 6656
rect 8205 6647 8263 6653
rect 8205 6613 8217 6647
rect 8251 6644 8263 6647
rect 10042 6644 10048 6656
rect 8251 6616 10048 6644
rect 8251 6613 8263 6616
rect 8205 6607 8263 6613
rect 10042 6604 10048 6616
rect 10100 6604 10106 6656
rect 12710 6604 12716 6656
rect 12768 6644 12774 6656
rect 13725 6647 13783 6653
rect 13725 6644 13737 6647
rect 12768 6616 13737 6644
rect 12768 6604 12774 6616
rect 13725 6613 13737 6616
rect 13771 6644 13783 6647
rect 16114 6644 16120 6656
rect 13771 6616 16120 6644
rect 13771 6613 13783 6616
rect 13725 6607 13783 6613
rect 16114 6604 16120 6616
rect 16172 6644 16178 6656
rect 16298 6644 16304 6656
rect 16172 6616 16304 6644
rect 16172 6604 16178 6616
rect 16298 6604 16304 6616
rect 16356 6604 16362 6656
rect 1104 6554 17388 6576
rect 1104 6502 3645 6554
rect 3697 6502 3709 6554
rect 3761 6502 3773 6554
rect 3825 6502 3837 6554
rect 3889 6502 3901 6554
rect 3953 6502 7716 6554
rect 7768 6502 7780 6554
rect 7832 6502 7844 6554
rect 7896 6502 7908 6554
rect 7960 6502 7972 6554
rect 8024 6502 11787 6554
rect 11839 6502 11851 6554
rect 11903 6502 11915 6554
rect 11967 6502 11979 6554
rect 12031 6502 12043 6554
rect 12095 6502 15858 6554
rect 15910 6502 15922 6554
rect 15974 6502 15986 6554
rect 16038 6502 16050 6554
rect 16102 6502 16114 6554
rect 16166 6502 17388 6554
rect 1104 6480 17388 6502
rect 2774 6400 2780 6452
rect 2832 6440 2838 6452
rect 3145 6443 3203 6449
rect 3145 6440 3157 6443
rect 2832 6412 3157 6440
rect 2832 6400 2838 6412
rect 3145 6409 3157 6412
rect 3191 6440 3203 6443
rect 5074 6440 5080 6452
rect 3191 6412 5080 6440
rect 3191 6409 3203 6412
rect 3145 6403 3203 6409
rect 5074 6400 5080 6412
rect 5132 6400 5138 6452
rect 6454 6400 6460 6452
rect 6512 6440 6518 6452
rect 11885 6443 11943 6449
rect 11885 6440 11897 6443
rect 6512 6412 11897 6440
rect 6512 6400 6518 6412
rect 11885 6409 11897 6412
rect 11931 6440 11943 6443
rect 14458 6440 14464 6452
rect 11931 6412 14464 6440
rect 11931 6409 11943 6412
rect 11885 6403 11943 6409
rect 14458 6400 14464 6412
rect 14516 6400 14522 6452
rect 9950 6332 9956 6384
rect 10008 6332 10014 6384
rect 10962 6332 10968 6384
rect 11020 6332 11026 6384
rect 11149 6375 11207 6381
rect 11149 6341 11161 6375
rect 11195 6372 11207 6375
rect 11195 6344 12020 6372
rect 11195 6341 11207 6344
rect 11149 6335 11207 6341
rect 2498 6264 2504 6316
rect 2556 6304 2562 6316
rect 3053 6307 3111 6313
rect 3053 6304 3065 6307
rect 2556 6276 3065 6304
rect 2556 6264 2562 6276
rect 3053 6273 3065 6276
rect 3099 6273 3111 6307
rect 3053 6267 3111 6273
rect 3329 6307 3387 6313
rect 3329 6273 3341 6307
rect 3375 6273 3387 6307
rect 3329 6267 3387 6273
rect 2866 6196 2872 6248
rect 2924 6236 2930 6248
rect 3344 6236 3372 6267
rect 8202 6264 8208 6316
rect 8260 6304 8266 6316
rect 8665 6307 8723 6313
rect 8665 6304 8677 6307
rect 8260 6276 8677 6304
rect 8260 6264 8266 6276
rect 8665 6273 8677 6276
rect 8711 6273 8723 6307
rect 8665 6267 8723 6273
rect 9122 6264 9128 6316
rect 9180 6304 9186 6316
rect 9217 6307 9275 6313
rect 9217 6304 9229 6307
rect 9180 6276 9229 6304
rect 9180 6264 9186 6276
rect 9217 6273 9229 6276
rect 9263 6273 9275 6307
rect 10980 6304 11008 6332
rect 11992 6313 12020 6344
rect 11057 6307 11115 6313
rect 11057 6304 11069 6307
rect 10980 6276 11069 6304
rect 9217 6267 9275 6273
rect 11057 6273 11069 6276
rect 11103 6273 11115 6307
rect 11057 6267 11115 6273
rect 11333 6307 11391 6313
rect 11333 6273 11345 6307
rect 11379 6304 11391 6307
rect 11701 6307 11759 6313
rect 11701 6304 11713 6307
rect 11379 6276 11713 6304
rect 11379 6273 11391 6276
rect 11333 6267 11391 6273
rect 11701 6273 11713 6276
rect 11747 6273 11759 6307
rect 11701 6267 11759 6273
rect 11977 6307 12035 6313
rect 11977 6273 11989 6307
rect 12023 6273 12035 6307
rect 11977 6267 12035 6273
rect 2924 6208 3372 6236
rect 9493 6239 9551 6245
rect 2924 6196 2930 6208
rect 9493 6205 9505 6239
rect 9539 6236 9551 6239
rect 9858 6236 9864 6248
rect 9539 6208 9864 6236
rect 9539 6205 9551 6208
rect 9493 6199 9551 6205
rect 9858 6196 9864 6208
rect 9916 6196 9922 6248
rect 10965 6239 11023 6245
rect 10965 6205 10977 6239
rect 11011 6236 11023 6239
rect 11348 6236 11376 6267
rect 11992 6236 12020 6267
rect 13722 6264 13728 6316
rect 13780 6264 13786 6316
rect 13817 6307 13875 6313
rect 13817 6273 13829 6307
rect 13863 6273 13875 6307
rect 13817 6267 13875 6273
rect 11011 6208 11376 6236
rect 11716 6208 12020 6236
rect 13832 6236 13860 6267
rect 13906 6264 13912 6316
rect 13964 6304 13970 6316
rect 14001 6307 14059 6313
rect 14001 6304 14013 6307
rect 13964 6276 14013 6304
rect 13964 6264 13970 6276
rect 14001 6273 14013 6276
rect 14047 6273 14059 6307
rect 14001 6267 14059 6273
rect 15746 6264 15752 6316
rect 15804 6264 15810 6316
rect 15933 6307 15991 6313
rect 15933 6273 15945 6307
rect 15979 6304 15991 6307
rect 16206 6304 16212 6316
rect 15979 6276 16212 6304
rect 15979 6273 15991 6276
rect 15933 6267 15991 6273
rect 16206 6264 16212 6276
rect 16264 6264 16270 6316
rect 14550 6236 14556 6248
rect 13832 6208 14556 6236
rect 11011 6205 11023 6208
rect 10965 6199 11023 6205
rect 11716 6180 11744 6208
rect 14550 6196 14556 6208
rect 14608 6196 14614 6248
rect 10778 6128 10784 6180
rect 10836 6168 10842 6180
rect 11057 6171 11115 6177
rect 11057 6168 11069 6171
rect 10836 6140 11069 6168
rect 10836 6128 10842 6140
rect 11057 6137 11069 6140
rect 11103 6137 11115 6171
rect 11057 6131 11115 6137
rect 11698 6128 11704 6180
rect 11756 6128 11762 6180
rect 3326 6060 3332 6112
rect 3384 6100 3390 6112
rect 3513 6103 3571 6109
rect 3513 6100 3525 6103
rect 3384 6072 3525 6100
rect 3384 6060 3390 6072
rect 3513 6069 3525 6072
rect 3559 6069 3571 6103
rect 3513 6063 3571 6069
rect 8941 6103 8999 6109
rect 8941 6069 8953 6103
rect 8987 6100 8999 6103
rect 10042 6100 10048 6112
rect 8987 6072 10048 6100
rect 8987 6069 8999 6072
rect 8941 6063 8999 6069
rect 10042 6060 10048 6072
rect 10100 6060 10106 6112
rect 10594 6060 10600 6112
rect 10652 6100 10658 6112
rect 11517 6103 11575 6109
rect 11517 6100 11529 6103
rect 10652 6072 11529 6100
rect 10652 6060 10658 6072
rect 11517 6069 11529 6072
rect 11563 6069 11575 6103
rect 11517 6063 11575 6069
rect 13909 6103 13967 6109
rect 13909 6069 13921 6103
rect 13955 6100 13967 6103
rect 13998 6100 14004 6112
rect 13955 6072 14004 6100
rect 13955 6069 13967 6072
rect 13909 6063 13967 6069
rect 13998 6060 14004 6072
rect 14056 6060 14062 6112
rect 15746 6060 15752 6112
rect 15804 6100 15810 6112
rect 15841 6103 15899 6109
rect 15841 6100 15853 6103
rect 15804 6072 15853 6100
rect 15804 6060 15810 6072
rect 15841 6069 15853 6072
rect 15887 6069 15899 6103
rect 15841 6063 15899 6069
rect 1104 6010 17388 6032
rect 1104 5958 2985 6010
rect 3037 5958 3049 6010
rect 3101 5958 3113 6010
rect 3165 5958 3177 6010
rect 3229 5958 3241 6010
rect 3293 5958 7056 6010
rect 7108 5958 7120 6010
rect 7172 5958 7184 6010
rect 7236 5958 7248 6010
rect 7300 5958 7312 6010
rect 7364 5958 11127 6010
rect 11179 5958 11191 6010
rect 11243 5958 11255 6010
rect 11307 5958 11319 6010
rect 11371 5958 11383 6010
rect 11435 5958 15198 6010
rect 15250 5958 15262 6010
rect 15314 5958 15326 6010
rect 15378 5958 15390 6010
rect 15442 5958 15454 6010
rect 15506 5958 17388 6010
rect 1104 5936 17388 5958
rect 3142 5856 3148 5908
rect 3200 5896 3206 5908
rect 3510 5896 3516 5908
rect 3200 5868 3516 5896
rect 3200 5856 3206 5868
rect 3510 5856 3516 5868
rect 3568 5856 3574 5908
rect 6914 5856 6920 5908
rect 6972 5896 6978 5908
rect 7190 5896 7196 5908
rect 6972 5868 7196 5896
rect 6972 5856 6978 5868
rect 7190 5856 7196 5868
rect 7248 5896 7254 5908
rect 8202 5896 8208 5908
rect 7248 5868 8208 5896
rect 7248 5856 7254 5868
rect 8202 5856 8208 5868
rect 8260 5856 8266 5908
rect 9858 5856 9864 5908
rect 9916 5856 9922 5908
rect 9950 5856 9956 5908
rect 10008 5896 10014 5908
rect 12434 5896 12440 5908
rect 10008 5868 12440 5896
rect 10008 5856 10014 5868
rect 12434 5856 12440 5868
rect 12492 5856 12498 5908
rect 13906 5856 13912 5908
rect 13964 5856 13970 5908
rect 1581 5831 1639 5837
rect 1581 5797 1593 5831
rect 1627 5828 1639 5831
rect 2498 5828 2504 5840
rect 1627 5800 2504 5828
rect 1627 5797 1639 5800
rect 1581 5791 1639 5797
rect 2498 5788 2504 5800
rect 2556 5788 2562 5840
rect 2593 5831 2651 5837
rect 2593 5797 2605 5831
rect 2639 5828 2651 5831
rect 2639 5800 3464 5828
rect 2639 5797 2651 5800
rect 2593 5791 2651 5797
rect 3436 5772 3464 5800
rect 7006 5788 7012 5840
rect 7064 5828 7070 5840
rect 7377 5831 7435 5837
rect 7377 5828 7389 5831
rect 7064 5800 7389 5828
rect 7064 5788 7070 5800
rect 7377 5797 7389 5800
rect 7423 5797 7435 5831
rect 7377 5791 7435 5797
rect 9125 5831 9183 5837
rect 9125 5797 9137 5831
rect 9171 5828 9183 5831
rect 10686 5828 10692 5840
rect 9171 5800 10692 5828
rect 9171 5797 9183 5800
rect 9125 5791 9183 5797
rect 10686 5788 10692 5800
rect 10744 5828 10750 5840
rect 10962 5828 10968 5840
rect 10744 5800 10968 5828
rect 10744 5788 10750 5800
rect 10962 5788 10968 5800
rect 11020 5788 11026 5840
rect 2961 5763 3019 5769
rect 2961 5729 2973 5763
rect 3007 5760 3019 5763
rect 3326 5760 3332 5772
rect 3007 5732 3332 5760
rect 3007 5729 3019 5732
rect 2961 5723 3019 5729
rect 3326 5720 3332 5732
rect 3384 5720 3390 5772
rect 3418 5720 3424 5772
rect 3476 5720 3482 5772
rect 3510 5720 3516 5772
rect 3568 5760 3574 5772
rect 3881 5763 3939 5769
rect 3881 5760 3893 5763
rect 3568 5732 3893 5760
rect 3568 5720 3574 5732
rect 3881 5729 3893 5732
rect 3927 5729 3939 5763
rect 3881 5723 3939 5729
rect 6822 5720 6828 5772
rect 6880 5760 6886 5772
rect 10045 5763 10103 5769
rect 6880 5732 7420 5760
rect 6880 5720 6886 5732
rect 1394 5652 1400 5704
rect 1452 5652 1458 5704
rect 2406 5652 2412 5704
rect 2464 5652 2470 5704
rect 2498 5652 2504 5704
rect 2556 5652 2562 5704
rect 2774 5652 2780 5704
rect 2832 5692 2838 5704
rect 3053 5695 3111 5701
rect 3053 5692 3065 5695
rect 2832 5664 3065 5692
rect 2832 5652 2838 5664
rect 3053 5661 3065 5664
rect 3099 5692 3111 5695
rect 3973 5695 4031 5701
rect 3973 5692 3985 5695
rect 3099 5664 3985 5692
rect 3099 5661 3111 5664
rect 3053 5655 3111 5661
rect 3973 5661 3985 5664
rect 4019 5661 4031 5695
rect 3973 5655 4031 5661
rect 6914 5652 6920 5704
rect 6972 5652 6978 5704
rect 7116 5701 7144 5732
rect 7101 5695 7159 5701
rect 7101 5661 7113 5695
rect 7147 5661 7159 5695
rect 7101 5655 7159 5661
rect 7190 5652 7196 5704
rect 7248 5652 7254 5704
rect 7392 5692 7420 5732
rect 10045 5729 10057 5763
rect 10091 5760 10103 5763
rect 10505 5763 10563 5769
rect 10091 5732 10456 5760
rect 10091 5729 10103 5732
rect 10045 5723 10103 5729
rect 7561 5695 7619 5701
rect 7561 5692 7573 5695
rect 7392 5664 7573 5692
rect 7561 5661 7573 5664
rect 7607 5661 7619 5695
rect 7561 5655 7619 5661
rect 8202 5652 8208 5704
rect 8260 5692 8266 5704
rect 8941 5695 8999 5701
rect 8941 5692 8953 5695
rect 8260 5664 8953 5692
rect 8260 5652 8266 5664
rect 8941 5661 8953 5664
rect 8987 5661 8999 5695
rect 8941 5655 8999 5661
rect 10134 5652 10140 5704
rect 10192 5652 10198 5704
rect 10428 5692 10456 5732
rect 10505 5729 10517 5763
rect 10551 5760 10563 5763
rect 10551 5732 10824 5760
rect 10551 5729 10563 5732
rect 10505 5723 10563 5729
rect 10796 5704 10824 5732
rect 11514 5720 11520 5772
rect 11572 5760 11578 5772
rect 12161 5763 12219 5769
rect 12161 5760 12173 5763
rect 11572 5732 12173 5760
rect 11572 5720 11578 5732
rect 12161 5729 12173 5732
rect 12207 5729 12219 5763
rect 12161 5723 12219 5729
rect 10594 5692 10600 5704
rect 10428 5664 10600 5692
rect 10594 5652 10600 5664
rect 10652 5652 10658 5704
rect 10778 5652 10784 5704
rect 10836 5652 10842 5704
rect 13924 5692 13952 5856
rect 14550 5788 14556 5840
rect 14608 5828 14614 5840
rect 16853 5831 16911 5837
rect 16853 5828 16865 5831
rect 14608 5800 16865 5828
rect 14608 5788 14614 5800
rect 16853 5797 16865 5800
rect 16899 5797 16911 5831
rect 16853 5791 16911 5797
rect 14277 5695 14335 5701
rect 14277 5692 14289 5695
rect 13924 5664 14289 5692
rect 14277 5661 14289 5664
rect 14323 5661 14335 5695
rect 14277 5655 14335 5661
rect 14458 5652 14464 5704
rect 14516 5652 14522 5704
rect 14568 5701 14596 5788
rect 15746 5720 15752 5772
rect 15804 5720 15810 5772
rect 14553 5695 14611 5701
rect 14553 5661 14565 5695
rect 14599 5661 14611 5695
rect 14553 5655 14611 5661
rect 15654 5652 15660 5704
rect 15712 5652 15718 5704
rect 17034 5652 17040 5704
rect 17092 5652 17098 5704
rect 2685 5627 2743 5633
rect 2685 5593 2697 5627
rect 2731 5624 2743 5627
rect 2866 5624 2872 5636
rect 2731 5596 2872 5624
rect 2731 5593 2743 5596
rect 2685 5587 2743 5593
rect 2866 5584 2872 5596
rect 2924 5624 2930 5636
rect 3234 5624 3240 5636
rect 2924 5596 3240 5624
rect 2924 5584 2930 5596
rect 3234 5584 3240 5596
rect 3292 5584 3298 5636
rect 5074 5584 5080 5636
rect 5132 5624 5138 5636
rect 6932 5624 6960 5652
rect 7285 5627 7343 5633
rect 7285 5624 7297 5627
rect 5132 5596 6868 5624
rect 6932 5596 7297 5624
rect 5132 5584 5138 5596
rect 2774 5516 2780 5568
rect 2832 5516 2838 5568
rect 4341 5559 4399 5565
rect 4341 5525 4353 5559
rect 4387 5556 4399 5559
rect 4522 5556 4528 5568
rect 4387 5528 4528 5556
rect 4387 5525 4399 5528
rect 4341 5519 4399 5525
rect 4522 5516 4528 5528
rect 4580 5516 4586 5568
rect 6546 5516 6552 5568
rect 6604 5556 6610 5568
rect 6733 5559 6791 5565
rect 6733 5556 6745 5559
rect 6604 5528 6745 5556
rect 6604 5516 6610 5528
rect 6733 5525 6745 5528
rect 6779 5525 6791 5559
rect 6840 5556 6868 5596
rect 7285 5593 7297 5596
rect 7331 5593 7343 5627
rect 7285 5587 7343 5593
rect 7469 5627 7527 5633
rect 7469 5593 7481 5627
rect 7515 5593 7527 5627
rect 7469 5587 7527 5593
rect 7484 5556 7512 5587
rect 12434 5584 12440 5636
rect 12492 5584 12498 5636
rect 12526 5584 12532 5636
rect 12584 5624 12590 5636
rect 12894 5624 12900 5636
rect 12584 5596 12900 5624
rect 12584 5584 12590 5596
rect 12894 5584 12900 5596
rect 12952 5584 12958 5636
rect 6840 5528 7512 5556
rect 6733 5519 6791 5525
rect 10594 5516 10600 5568
rect 10652 5516 10658 5568
rect 14090 5516 14096 5568
rect 14148 5516 14154 5568
rect 16025 5559 16083 5565
rect 16025 5525 16037 5559
rect 16071 5556 16083 5559
rect 16758 5556 16764 5568
rect 16071 5528 16764 5556
rect 16071 5525 16083 5528
rect 16025 5519 16083 5525
rect 16758 5516 16764 5528
rect 16816 5516 16822 5568
rect 1104 5466 17388 5488
rect 1104 5414 3645 5466
rect 3697 5414 3709 5466
rect 3761 5414 3773 5466
rect 3825 5414 3837 5466
rect 3889 5414 3901 5466
rect 3953 5414 7716 5466
rect 7768 5414 7780 5466
rect 7832 5414 7844 5466
rect 7896 5414 7908 5466
rect 7960 5414 7972 5466
rect 8024 5414 11787 5466
rect 11839 5414 11851 5466
rect 11903 5414 11915 5466
rect 11967 5414 11979 5466
rect 12031 5414 12043 5466
rect 12095 5414 15858 5466
rect 15910 5414 15922 5466
rect 15974 5414 15986 5466
rect 16038 5414 16050 5466
rect 16102 5414 16114 5466
rect 16166 5414 17388 5466
rect 1104 5392 17388 5414
rect 2774 5352 2780 5364
rect 1872 5324 2780 5352
rect 1872 5293 1900 5324
rect 2774 5312 2780 5324
rect 2832 5312 2838 5364
rect 3510 5312 3516 5364
rect 3568 5312 3574 5364
rect 7006 5312 7012 5364
rect 7064 5352 7070 5364
rect 7374 5352 7380 5364
rect 7064 5324 7380 5352
rect 7064 5312 7070 5324
rect 7374 5312 7380 5324
rect 7432 5312 7438 5364
rect 7653 5355 7711 5361
rect 7653 5321 7665 5355
rect 7699 5321 7711 5355
rect 7653 5315 7711 5321
rect 1857 5287 1915 5293
rect 1857 5253 1869 5287
rect 1903 5253 1915 5287
rect 3142 5284 3148 5296
rect 3082 5256 3148 5284
rect 1857 5247 1915 5253
rect 3142 5244 3148 5256
rect 3200 5244 3206 5296
rect 3326 5244 3332 5296
rect 3384 5284 3390 5296
rect 3384 5256 3648 5284
rect 3384 5244 3390 5256
rect 3418 5176 3424 5228
rect 3476 5176 3482 5228
rect 3620 5225 3648 5256
rect 4522 5244 4528 5296
rect 4580 5244 4586 5296
rect 5258 5244 5264 5296
rect 5316 5244 5322 5296
rect 7668 5284 7696 5315
rect 7742 5312 7748 5364
rect 7800 5352 7806 5364
rect 9677 5355 9735 5361
rect 7800 5324 8340 5352
rect 7800 5312 7806 5324
rect 8205 5287 8263 5293
rect 8205 5284 8217 5287
rect 7668 5256 8217 5284
rect 8205 5253 8217 5256
rect 8251 5253 8263 5287
rect 8312 5284 8340 5324
rect 9677 5321 9689 5355
rect 9723 5352 9735 5355
rect 10134 5352 10140 5364
rect 9723 5324 10140 5352
rect 9723 5321 9735 5324
rect 9677 5315 9735 5321
rect 10134 5312 10140 5324
rect 10192 5312 10198 5364
rect 10873 5355 10931 5361
rect 10873 5321 10885 5355
rect 10919 5321 10931 5355
rect 10873 5315 10931 5321
rect 8312 5256 8694 5284
rect 8205 5247 8263 5253
rect 3605 5219 3663 5225
rect 3605 5185 3617 5219
rect 3651 5185 3663 5219
rect 7285 5219 7343 5225
rect 7285 5216 7297 5219
rect 3605 5179 3663 5185
rect 6656 5188 7297 5216
rect 1578 5108 1584 5160
rect 1636 5108 1642 5160
rect 4154 5148 4160 5160
rect 3252 5120 4160 5148
rect 1596 5012 1624 5108
rect 3252 5012 3280 5120
rect 4154 5108 4160 5120
rect 4212 5148 4218 5160
rect 4249 5151 4307 5157
rect 4249 5148 4261 5151
rect 4212 5120 4261 5148
rect 4212 5108 4218 5120
rect 4249 5117 4261 5120
rect 4295 5148 4307 5151
rect 5074 5148 5080 5160
rect 4295 5120 5080 5148
rect 4295 5117 4307 5120
rect 4249 5111 4307 5117
rect 5074 5108 5080 5120
rect 5132 5108 5138 5160
rect 6546 5108 6552 5160
rect 6604 5108 6610 5160
rect 6656 5157 6684 5188
rect 7285 5185 7297 5188
rect 7331 5185 7343 5219
rect 10152 5216 10180 5312
rect 10888 5284 10916 5315
rect 12434 5312 12440 5364
rect 12492 5352 12498 5364
rect 13357 5355 13415 5361
rect 13357 5352 13369 5355
rect 12492 5324 13369 5352
rect 12492 5312 12498 5324
rect 13357 5321 13369 5324
rect 13403 5321 13415 5355
rect 13357 5315 13415 5321
rect 13998 5312 14004 5364
rect 14056 5312 14062 5364
rect 15562 5312 15568 5364
rect 15620 5352 15626 5364
rect 16025 5355 16083 5361
rect 16025 5352 16037 5355
rect 15620 5324 16037 5352
rect 15620 5312 15626 5324
rect 16025 5321 16037 5324
rect 16071 5321 16083 5355
rect 16025 5315 16083 5321
rect 11793 5287 11851 5293
rect 11793 5284 11805 5287
rect 10888 5256 11805 5284
rect 11793 5253 11805 5256
rect 11839 5253 11851 5287
rect 11793 5247 11851 5253
rect 12526 5244 12532 5296
rect 12584 5244 12590 5296
rect 14458 5284 14464 5296
rect 14292 5256 14464 5284
rect 10505 5219 10563 5225
rect 10505 5216 10517 5219
rect 10152 5188 10517 5216
rect 7285 5179 7343 5185
rect 10505 5185 10517 5188
rect 10551 5185 10563 5219
rect 10505 5179 10563 5185
rect 11514 5176 11520 5228
rect 11572 5176 11578 5228
rect 13541 5219 13599 5225
rect 13541 5185 13553 5219
rect 13587 5216 13599 5219
rect 14090 5216 14096 5228
rect 13587 5188 14096 5216
rect 13587 5185 13599 5188
rect 13541 5179 13599 5185
rect 14090 5176 14096 5188
rect 14148 5176 14154 5228
rect 14292 5225 14320 5256
rect 14458 5244 14464 5256
rect 14516 5284 14522 5296
rect 14642 5284 14648 5296
rect 14516 5256 14648 5284
rect 14516 5244 14522 5256
rect 14642 5244 14648 5256
rect 14700 5244 14706 5296
rect 14277 5219 14335 5225
rect 14277 5185 14289 5219
rect 14323 5185 14335 5219
rect 16390 5216 16396 5228
rect 15686 5188 16396 5216
rect 14277 5179 14335 5185
rect 15764 5160 15792 5188
rect 16390 5176 16396 5188
rect 16448 5176 16454 5228
rect 6641 5151 6699 5157
rect 6641 5117 6653 5151
rect 6687 5117 6699 5151
rect 6641 5111 6699 5117
rect 7377 5151 7435 5157
rect 7377 5117 7389 5151
rect 7423 5148 7435 5151
rect 7558 5148 7564 5160
rect 7423 5120 7564 5148
rect 7423 5117 7435 5120
rect 7377 5111 7435 5117
rect 3326 5040 3332 5092
rect 3384 5040 3390 5092
rect 5997 5083 6055 5089
rect 5997 5049 6009 5083
rect 6043 5080 6055 5083
rect 6656 5080 6684 5111
rect 7558 5108 7564 5120
rect 7616 5108 7622 5160
rect 7929 5151 7987 5157
rect 7929 5117 7941 5151
rect 7975 5148 7987 5151
rect 8202 5148 8208 5160
rect 7975 5120 8208 5148
rect 7975 5117 7987 5120
rect 7929 5111 7987 5117
rect 6043 5052 6684 5080
rect 6043 5049 6055 5052
rect 5997 5043 6055 5049
rect 7282 5040 7288 5092
rect 7340 5080 7346 5092
rect 7944 5080 7972 5111
rect 8202 5108 8208 5120
rect 8260 5108 8266 5160
rect 10594 5108 10600 5160
rect 10652 5108 10658 5160
rect 13633 5151 13691 5157
rect 13633 5117 13645 5151
rect 13679 5117 13691 5151
rect 13633 5111 13691 5117
rect 7340 5052 7972 5080
rect 13265 5083 13323 5089
rect 7340 5040 7346 5052
rect 13265 5049 13277 5083
rect 13311 5080 13323 5083
rect 13648 5080 13676 5111
rect 14550 5108 14556 5160
rect 14608 5108 14614 5160
rect 15746 5108 15752 5160
rect 15804 5108 15810 5160
rect 13311 5052 14320 5080
rect 13311 5049 13323 5052
rect 13265 5043 13323 5049
rect 14292 5024 14320 5052
rect 1596 4984 3280 5012
rect 6362 4972 6368 5024
rect 6420 4972 6426 5024
rect 14274 4972 14280 5024
rect 14332 4972 14338 5024
rect 1104 4922 17388 4944
rect 1104 4870 2985 4922
rect 3037 4870 3049 4922
rect 3101 4870 3113 4922
rect 3165 4870 3177 4922
rect 3229 4870 3241 4922
rect 3293 4870 7056 4922
rect 7108 4870 7120 4922
rect 7172 4870 7184 4922
rect 7236 4870 7248 4922
rect 7300 4870 7312 4922
rect 7364 4870 11127 4922
rect 11179 4870 11191 4922
rect 11243 4870 11255 4922
rect 11307 4870 11319 4922
rect 11371 4870 11383 4922
rect 11435 4870 15198 4922
rect 15250 4870 15262 4922
rect 15314 4870 15326 4922
rect 15378 4870 15390 4922
rect 15442 4870 15454 4922
rect 15506 4870 17388 4922
rect 1104 4848 17388 4870
rect 6825 4811 6883 4817
rect 6825 4777 6837 4811
rect 6871 4808 6883 4811
rect 6914 4808 6920 4820
rect 6871 4780 6920 4808
rect 6871 4777 6883 4780
rect 6825 4771 6883 4777
rect 6914 4768 6920 4780
rect 6972 4768 6978 4820
rect 7558 4768 7564 4820
rect 7616 4768 7622 4820
rect 14550 4768 14556 4820
rect 14608 4768 14614 4820
rect 15764 4780 16988 4808
rect 14090 4740 14096 4752
rect 13556 4712 14096 4740
rect 5074 4632 5080 4684
rect 5132 4632 5138 4684
rect 5353 4675 5411 4681
rect 5353 4641 5365 4675
rect 5399 4672 5411 4675
rect 6362 4672 6368 4684
rect 5399 4644 6368 4672
rect 5399 4641 5411 4644
rect 5353 4635 5411 4641
rect 6362 4632 6368 4644
rect 6420 4632 6426 4684
rect 6546 4632 6552 4684
rect 6604 4632 6610 4684
rect 7374 4632 7380 4684
rect 7432 4672 7438 4684
rect 7432 4644 7696 4672
rect 7432 4632 7438 4644
rect 6564 4604 6592 4632
rect 7668 4613 7696 4644
rect 13556 4613 13584 4712
rect 14090 4700 14096 4712
rect 14148 4700 14154 4752
rect 14458 4700 14464 4752
rect 14516 4740 14522 4752
rect 15764 4740 15792 4780
rect 14516 4712 15792 4740
rect 14516 4700 14522 4712
rect 13633 4675 13691 4681
rect 13633 4641 13645 4675
rect 13679 4672 13691 4675
rect 14185 4675 14243 4681
rect 14185 4672 14197 4675
rect 13679 4644 14197 4672
rect 13679 4641 13691 4644
rect 13633 4635 13691 4641
rect 14185 4641 14197 4644
rect 14231 4641 14243 4675
rect 14185 4635 14243 4641
rect 16758 4632 16764 4684
rect 16816 4632 16822 4684
rect 16960 4672 16988 4780
rect 17037 4675 17095 4681
rect 17037 4672 17049 4675
rect 16960 4644 17049 4672
rect 17037 4641 17049 4644
rect 17083 4641 17095 4675
rect 17037 4635 17095 4641
rect 7469 4607 7527 4613
rect 7469 4604 7481 4607
rect 6564 4576 7481 4604
rect 7469 4573 7481 4576
rect 7515 4573 7527 4607
rect 7469 4567 7527 4573
rect 7653 4607 7711 4613
rect 7653 4573 7665 4607
rect 7699 4573 7711 4607
rect 7653 4567 7711 4573
rect 13541 4607 13599 4613
rect 13541 4573 13553 4607
rect 13587 4573 13599 4607
rect 13541 4567 13599 4573
rect 13725 4607 13783 4613
rect 13725 4573 13737 4607
rect 13771 4604 13783 4607
rect 13998 4604 14004 4616
rect 13771 4576 14004 4604
rect 13771 4573 13783 4576
rect 13725 4567 13783 4573
rect 13998 4564 14004 4576
rect 14056 4564 14062 4616
rect 14274 4564 14280 4616
rect 14332 4564 14338 4616
rect 6917 4539 6975 4545
rect 6917 4536 6929 4539
rect 6578 4508 6929 4536
rect 5258 4428 5264 4480
rect 5316 4468 5322 4480
rect 6656 4468 6684 4508
rect 6917 4505 6929 4508
rect 6963 4505 6975 4539
rect 6917 4499 6975 4505
rect 7285 4539 7343 4545
rect 7285 4505 7297 4539
rect 7331 4536 7343 4539
rect 10226 4536 10232 4548
rect 7331 4508 10232 4536
rect 7331 4505 7343 4508
rect 7285 4499 7343 4505
rect 10226 4496 10232 4508
rect 10284 4496 10290 4548
rect 15746 4496 15752 4548
rect 15804 4496 15810 4548
rect 5316 4440 6684 4468
rect 5316 4428 5322 4440
rect 15286 4428 15292 4480
rect 15344 4428 15350 4480
rect 1104 4378 17388 4400
rect 1104 4326 3645 4378
rect 3697 4326 3709 4378
rect 3761 4326 3773 4378
rect 3825 4326 3837 4378
rect 3889 4326 3901 4378
rect 3953 4326 7716 4378
rect 7768 4326 7780 4378
rect 7832 4326 7844 4378
rect 7896 4326 7908 4378
rect 7960 4326 7972 4378
rect 8024 4326 11787 4378
rect 11839 4326 11851 4378
rect 11903 4326 11915 4378
rect 11967 4326 11979 4378
rect 12031 4326 12043 4378
rect 12095 4326 15858 4378
rect 15910 4326 15922 4378
rect 15974 4326 15986 4378
rect 16038 4326 16050 4378
rect 16102 4326 16114 4378
rect 16166 4326 17388 4378
rect 1104 4304 17388 4326
rect 5166 4224 5172 4276
rect 5224 4264 5230 4276
rect 5261 4267 5319 4273
rect 5261 4264 5273 4267
rect 5224 4236 5273 4264
rect 5224 4224 5230 4236
rect 5261 4233 5273 4236
rect 5307 4264 5319 4267
rect 5810 4264 5816 4276
rect 5307 4236 5816 4264
rect 5307 4233 5319 4236
rect 5261 4227 5319 4233
rect 5810 4224 5816 4236
rect 5868 4224 5874 4276
rect 8864 4236 9628 4264
rect 7558 4156 7564 4208
rect 7616 4196 7622 4208
rect 8864 4196 8892 4236
rect 7616 4168 8970 4196
rect 7616 4156 7622 4168
rect 5074 4088 5080 4140
rect 5132 4088 5138 4140
rect 5353 4131 5411 4137
rect 5353 4097 5365 4131
rect 5399 4128 5411 4131
rect 5442 4128 5448 4140
rect 5399 4100 5448 4128
rect 5399 4097 5411 4100
rect 5353 4091 5411 4097
rect 5442 4088 5448 4100
rect 5500 4088 5506 4140
rect 8202 4088 8208 4140
rect 8260 4088 8266 4140
rect 9600 4128 9628 4236
rect 10226 4156 10232 4208
rect 10284 4196 10290 4208
rect 12986 4196 12992 4208
rect 10284 4168 12992 4196
rect 10284 4156 10290 4168
rect 12986 4156 12992 4168
rect 13044 4196 13050 4208
rect 13044 4168 13768 4196
rect 13044 4156 13050 4168
rect 10045 4131 10103 4137
rect 10045 4128 10057 4131
rect 9600 4114 10057 4128
rect 9614 4100 10057 4114
rect 10045 4097 10057 4100
rect 10091 4097 10103 4131
rect 10045 4091 10103 4097
rect 12529 4131 12587 4137
rect 12529 4097 12541 4131
rect 12575 4128 12587 4131
rect 12618 4128 12624 4140
rect 12575 4100 12624 4128
rect 12575 4097 12587 4100
rect 12529 4091 12587 4097
rect 12618 4088 12624 4100
rect 12676 4088 12682 4140
rect 12710 4088 12716 4140
rect 12768 4088 12774 4140
rect 12805 4131 12863 4137
rect 12805 4097 12817 4131
rect 12851 4128 12863 4131
rect 13446 4128 13452 4140
rect 12851 4100 13452 4128
rect 12851 4097 12863 4100
rect 12805 4091 12863 4097
rect 13446 4088 13452 4100
rect 13504 4088 13510 4140
rect 8481 4063 8539 4069
rect 8481 4029 8493 4063
rect 8527 4060 8539 4063
rect 8938 4060 8944 4072
rect 8527 4032 8944 4060
rect 8527 4029 8539 4032
rect 8481 4023 8539 4029
rect 8938 4020 8944 4032
rect 8996 4020 9002 4072
rect 10042 3952 10048 4004
rect 10100 3992 10106 4004
rect 12728 3992 12756 4088
rect 10100 3964 12756 3992
rect 13740 3992 13768 4168
rect 14921 4131 14979 4137
rect 14921 4097 14933 4131
rect 14967 4128 14979 4131
rect 15286 4128 15292 4140
rect 14967 4100 15292 4128
rect 14967 4097 14979 4100
rect 14921 4091 14979 4097
rect 15286 4088 15292 4100
rect 15344 4088 15350 4140
rect 15470 4088 15476 4140
rect 15528 4088 15534 4140
rect 15562 4088 15568 4140
rect 15620 4088 15626 4140
rect 15749 4131 15807 4137
rect 15749 4097 15761 4131
rect 15795 4128 15807 4131
rect 16574 4128 16580 4140
rect 15795 4100 16580 4128
rect 15795 4097 15807 4100
rect 15749 4091 15807 4097
rect 16574 4088 16580 4100
rect 16632 4088 16638 4140
rect 15013 4063 15071 4069
rect 15013 4029 15025 4063
rect 15059 4060 15071 4063
rect 15657 4063 15715 4069
rect 15657 4060 15669 4063
rect 15059 4032 15669 4060
rect 15059 4029 15071 4032
rect 15013 4023 15071 4029
rect 15657 4029 15669 4032
rect 15703 4029 15715 4063
rect 15657 4023 15715 4029
rect 15289 3995 15347 4001
rect 15289 3992 15301 3995
rect 13740 3964 15301 3992
rect 10100 3952 10106 3964
rect 15289 3961 15301 3964
rect 15335 3992 15347 3995
rect 16482 3992 16488 4004
rect 15335 3964 16488 3992
rect 15335 3961 15347 3964
rect 15289 3955 15347 3961
rect 15672 3936 15700 3964
rect 16482 3952 16488 3964
rect 16540 3952 16546 4004
rect 4706 3884 4712 3936
rect 4764 3924 4770 3936
rect 4893 3927 4951 3933
rect 4893 3924 4905 3927
rect 4764 3896 4905 3924
rect 4764 3884 4770 3896
rect 4893 3893 4905 3896
rect 4939 3893 4951 3927
rect 4893 3887 4951 3893
rect 9858 3884 9864 3936
rect 9916 3924 9922 3936
rect 9953 3927 10011 3933
rect 9953 3924 9965 3927
rect 9916 3896 9965 3924
rect 9916 3884 9922 3896
rect 9953 3893 9965 3896
rect 9999 3893 10011 3927
rect 9953 3887 10011 3893
rect 12250 3884 12256 3936
rect 12308 3924 12314 3936
rect 12345 3927 12403 3933
rect 12345 3924 12357 3927
rect 12308 3896 12357 3924
rect 12308 3884 12314 3896
rect 12345 3893 12357 3896
rect 12391 3893 12403 3927
rect 12345 3887 12403 3893
rect 14090 3884 14096 3936
rect 14148 3924 14154 3936
rect 14645 3927 14703 3933
rect 14645 3924 14657 3927
rect 14148 3896 14657 3924
rect 14148 3884 14154 3896
rect 14645 3893 14657 3896
rect 14691 3893 14703 3927
rect 14645 3887 14703 3893
rect 15654 3884 15660 3936
rect 15712 3884 15718 3936
rect 1104 3834 17388 3856
rect 1104 3782 2985 3834
rect 3037 3782 3049 3834
rect 3101 3782 3113 3834
rect 3165 3782 3177 3834
rect 3229 3782 3241 3834
rect 3293 3782 7056 3834
rect 7108 3782 7120 3834
rect 7172 3782 7184 3834
rect 7236 3782 7248 3834
rect 7300 3782 7312 3834
rect 7364 3782 11127 3834
rect 11179 3782 11191 3834
rect 11243 3782 11255 3834
rect 11307 3782 11319 3834
rect 11371 3782 11383 3834
rect 11435 3782 15198 3834
rect 15250 3782 15262 3834
rect 15314 3782 15326 3834
rect 15378 3782 15390 3834
rect 15442 3782 15454 3834
rect 15506 3782 17388 3834
rect 1104 3760 17388 3782
rect 5074 3680 5080 3732
rect 5132 3720 5138 3732
rect 5537 3723 5595 3729
rect 5537 3720 5549 3723
rect 5132 3692 5549 3720
rect 5132 3680 5138 3692
rect 5537 3689 5549 3692
rect 5583 3689 5595 3723
rect 5537 3683 5595 3689
rect 7745 3723 7803 3729
rect 7745 3689 7757 3723
rect 7791 3720 7803 3723
rect 8110 3720 8116 3732
rect 7791 3692 8116 3720
rect 7791 3689 7803 3692
rect 7745 3683 7803 3689
rect 3789 3587 3847 3593
rect 3789 3553 3801 3587
rect 3835 3584 3847 3587
rect 4154 3584 4160 3596
rect 3835 3556 4160 3584
rect 3835 3553 3847 3556
rect 3789 3547 3847 3553
rect 4154 3544 4160 3556
rect 4212 3544 4218 3596
rect 5258 3584 5264 3596
rect 5184 3556 5264 3584
rect 5184 3502 5212 3556
rect 5258 3544 5264 3556
rect 5316 3544 5322 3596
rect 5552 3516 5580 3683
rect 8110 3680 8116 3692
rect 8168 3680 8174 3732
rect 8938 3680 8944 3732
rect 8996 3680 9002 3732
rect 12618 3680 12624 3732
rect 12676 3680 12682 3732
rect 12894 3680 12900 3732
rect 12952 3680 12958 3732
rect 13722 3720 13728 3732
rect 13556 3692 13728 3720
rect 10321 3655 10379 3661
rect 10321 3621 10333 3655
rect 10367 3621 10379 3655
rect 10321 3615 10379 3621
rect 5997 3587 6055 3593
rect 5997 3553 6009 3587
rect 6043 3584 6055 3587
rect 8202 3584 8208 3596
rect 6043 3556 8208 3584
rect 6043 3553 6055 3556
rect 5997 3547 6055 3553
rect 8202 3544 8208 3556
rect 8260 3544 8266 3596
rect 9125 3587 9183 3593
rect 9125 3584 9137 3587
rect 8588 3556 9137 3584
rect 8588 3525 8616 3556
rect 9125 3553 9137 3556
rect 9171 3584 9183 3587
rect 9677 3587 9735 3593
rect 9677 3584 9689 3587
rect 9171 3556 9689 3584
rect 9171 3553 9183 3556
rect 9125 3547 9183 3553
rect 9677 3553 9689 3556
rect 9723 3553 9735 3587
rect 10336 3584 10364 3615
rect 9677 3547 9735 3553
rect 9784 3556 10364 3584
rect 10873 3587 10931 3593
rect 5905 3519 5963 3525
rect 5905 3516 5917 3519
rect 5552 3488 5917 3516
rect 5905 3485 5917 3488
rect 5951 3485 5963 3519
rect 5905 3479 5963 3485
rect 8573 3519 8631 3525
rect 8573 3485 8585 3519
rect 8619 3485 8631 3519
rect 8573 3479 8631 3485
rect 8757 3519 8815 3525
rect 8757 3485 8769 3519
rect 8803 3485 8815 3519
rect 8757 3479 8815 3485
rect 4062 3408 4068 3460
rect 4120 3408 4126 3460
rect 5442 3408 5448 3460
rect 5500 3448 5506 3460
rect 5629 3451 5687 3457
rect 5629 3448 5641 3451
rect 5500 3420 5641 3448
rect 5500 3408 5506 3420
rect 5629 3417 5641 3420
rect 5675 3417 5687 3451
rect 5629 3411 5687 3417
rect 5810 3408 5816 3460
rect 5868 3408 5874 3460
rect 6270 3408 6276 3460
rect 6328 3408 6334 3460
rect 7558 3448 7564 3460
rect 7498 3420 7564 3448
rect 7558 3408 7564 3420
rect 7616 3408 7622 3460
rect 8772 3448 8800 3479
rect 9030 3476 9036 3528
rect 9088 3516 9094 3528
rect 9217 3519 9275 3525
rect 9217 3516 9229 3519
rect 9088 3488 9229 3516
rect 9088 3476 9094 3488
rect 9217 3485 9229 3488
rect 9263 3485 9275 3519
rect 9217 3479 9275 3485
rect 9585 3519 9643 3525
rect 9585 3485 9597 3519
rect 9631 3516 9643 3519
rect 9784 3516 9812 3556
rect 10873 3553 10885 3587
rect 10919 3584 10931 3587
rect 11514 3584 11520 3596
rect 10919 3556 11520 3584
rect 10919 3553 10931 3556
rect 10873 3547 10931 3553
rect 11514 3544 11520 3556
rect 11572 3544 11578 3596
rect 9631 3488 9812 3516
rect 9631 3485 9643 3488
rect 9585 3479 9643 3485
rect 9600 3448 9628 3479
rect 9858 3476 9864 3528
rect 9916 3476 9922 3528
rect 10042 3476 10048 3528
rect 10100 3476 10106 3528
rect 10134 3476 10140 3528
rect 10192 3516 10198 3528
rect 10413 3519 10471 3525
rect 10413 3516 10425 3519
rect 10192 3488 10425 3516
rect 10192 3476 10198 3488
rect 10413 3485 10425 3488
rect 10459 3485 10471 3519
rect 10413 3479 10471 3485
rect 10505 3519 10563 3525
rect 10505 3485 10517 3519
rect 10551 3516 10563 3519
rect 10686 3516 10692 3528
rect 10551 3488 10692 3516
rect 10551 3485 10563 3488
rect 10505 3479 10563 3485
rect 10686 3476 10692 3488
rect 10744 3476 10750 3528
rect 12636 3516 12664 3680
rect 13265 3519 13323 3525
rect 13265 3516 13277 3519
rect 12636 3488 13277 3516
rect 13265 3485 13277 3488
rect 13311 3485 13323 3519
rect 13265 3479 13323 3485
rect 13446 3476 13452 3528
rect 13504 3476 13510 3528
rect 13556 3525 13584 3692
rect 13722 3680 13728 3692
rect 13780 3720 13786 3732
rect 13780 3692 15424 3720
rect 13780 3680 13786 3692
rect 15396 3652 15424 3692
rect 16574 3680 16580 3732
rect 16632 3680 16638 3732
rect 16850 3652 16856 3664
rect 15396 3624 16856 3652
rect 14093 3587 14151 3593
rect 14093 3553 14105 3587
rect 14139 3584 14151 3587
rect 14458 3584 14464 3596
rect 14139 3556 14464 3584
rect 14139 3553 14151 3556
rect 14093 3547 14151 3553
rect 14458 3544 14464 3556
rect 14516 3544 14522 3596
rect 15841 3587 15899 3593
rect 15841 3553 15853 3587
rect 15887 3584 15899 3587
rect 15887 3556 16160 3584
rect 15887 3553 15899 3556
rect 15841 3547 15899 3553
rect 16132 3525 16160 3556
rect 13541 3519 13599 3525
rect 13541 3485 13553 3519
rect 13587 3485 13599 3519
rect 13541 3479 13599 3485
rect 16117 3519 16175 3525
rect 16117 3485 16129 3519
rect 16163 3485 16175 3519
rect 16117 3479 16175 3485
rect 8772 3420 9628 3448
rect 9876 3448 9904 3476
rect 10229 3451 10287 3457
rect 10229 3448 10241 3451
rect 9876 3420 10241 3448
rect 10229 3417 10241 3420
rect 10275 3417 10287 3451
rect 10229 3411 10287 3417
rect 11146 3408 11152 3460
rect 11204 3408 11210 3460
rect 11606 3448 11612 3460
rect 11532 3420 11612 3448
rect 5905 3383 5963 3389
rect 5905 3349 5917 3383
rect 5951 3380 5963 3383
rect 6086 3380 6092 3392
rect 5951 3352 6092 3380
rect 5951 3349 5963 3352
rect 5905 3343 5963 3349
rect 6086 3340 6092 3352
rect 6144 3340 6150 3392
rect 8662 3340 8668 3392
rect 8720 3340 8726 3392
rect 11532 3380 11560 3420
rect 11606 3408 11612 3420
rect 11664 3408 11670 3460
rect 12805 3451 12863 3457
rect 12805 3417 12817 3451
rect 12851 3448 12863 3451
rect 12986 3448 12992 3460
rect 12851 3420 12992 3448
rect 12851 3417 12863 3420
rect 12805 3411 12863 3417
rect 12986 3408 12992 3420
rect 13044 3408 13050 3460
rect 14369 3451 14427 3457
rect 14369 3417 14381 3451
rect 14415 3448 14427 3451
rect 14642 3448 14648 3460
rect 14415 3420 14648 3448
rect 14415 3417 14427 3420
rect 14369 3411 14427 3417
rect 14642 3408 14648 3420
rect 14700 3408 14706 3460
rect 15838 3448 15844 3460
rect 14752 3420 14858 3448
rect 15672 3420 15844 3448
rect 12894 3380 12900 3392
rect 11532 3352 12900 3380
rect 12894 3340 12900 3352
rect 12952 3340 12958 3392
rect 13354 3340 13360 3392
rect 13412 3340 13418 3392
rect 13630 3340 13636 3392
rect 13688 3380 13694 3392
rect 14752 3380 14780 3420
rect 15378 3380 15384 3392
rect 13688 3352 15384 3380
rect 13688 3340 13694 3352
rect 15378 3340 15384 3352
rect 15436 3380 15442 3392
rect 15672 3380 15700 3420
rect 15838 3408 15844 3420
rect 15896 3408 15902 3460
rect 16132 3448 16160 3479
rect 16298 3476 16304 3528
rect 16356 3476 16362 3528
rect 16776 3525 16804 3624
rect 16850 3612 16856 3624
rect 16908 3612 16914 3664
rect 16393 3519 16451 3525
rect 16393 3485 16405 3519
rect 16439 3516 16451 3519
rect 16761 3519 16819 3525
rect 16439 3488 16712 3516
rect 16439 3485 16451 3488
rect 16393 3479 16451 3485
rect 16684 3457 16712 3488
rect 16761 3485 16773 3519
rect 16807 3485 16819 3519
rect 16761 3479 16819 3485
rect 17034 3476 17040 3528
rect 17092 3476 17098 3528
rect 16485 3451 16543 3457
rect 16485 3448 16497 3451
rect 16132 3420 16497 3448
rect 16485 3417 16497 3420
rect 16531 3417 16543 3451
rect 16485 3411 16543 3417
rect 16669 3451 16727 3457
rect 16669 3417 16681 3451
rect 16715 3417 16727 3451
rect 16669 3411 16727 3417
rect 15436 3352 15700 3380
rect 15436 3340 15442 3352
rect 15746 3340 15752 3392
rect 15804 3380 15810 3392
rect 15933 3383 15991 3389
rect 15933 3380 15945 3383
rect 15804 3352 15945 3380
rect 15804 3340 15810 3352
rect 15933 3349 15945 3352
rect 15979 3349 15991 3383
rect 16684 3380 16712 3411
rect 16853 3383 16911 3389
rect 16853 3380 16865 3383
rect 16684 3352 16865 3380
rect 15933 3343 15991 3349
rect 16853 3349 16865 3352
rect 16899 3349 16911 3383
rect 16853 3343 16911 3349
rect 1104 3290 17388 3312
rect 1104 3238 3645 3290
rect 3697 3238 3709 3290
rect 3761 3238 3773 3290
rect 3825 3238 3837 3290
rect 3889 3238 3901 3290
rect 3953 3238 7716 3290
rect 7768 3238 7780 3290
rect 7832 3238 7844 3290
rect 7896 3238 7908 3290
rect 7960 3238 7972 3290
rect 8024 3238 11787 3290
rect 11839 3238 11851 3290
rect 11903 3238 11915 3290
rect 11967 3238 11979 3290
rect 12031 3238 12043 3290
rect 12095 3238 15858 3290
rect 15910 3238 15922 3290
rect 15974 3238 15986 3290
rect 16038 3238 16050 3290
rect 16102 3238 16114 3290
rect 16166 3238 17388 3290
rect 1104 3216 17388 3238
rect 4062 3136 4068 3188
rect 4120 3176 4126 3188
rect 4525 3179 4583 3185
rect 4525 3176 4537 3179
rect 4120 3148 4537 3176
rect 4120 3136 4126 3148
rect 4525 3145 4537 3148
rect 4571 3145 4583 3179
rect 4525 3139 4583 3145
rect 4706 3136 4712 3188
rect 4764 3176 4770 3188
rect 5718 3176 5724 3188
rect 4764 3148 5724 3176
rect 4764 3136 4770 3148
rect 5718 3136 5724 3148
rect 5776 3136 5782 3188
rect 5813 3179 5871 3185
rect 5813 3145 5825 3179
rect 5859 3176 5871 3179
rect 6270 3176 6276 3188
rect 5859 3148 6276 3176
rect 5859 3145 5871 3148
rect 5813 3139 5871 3145
rect 6270 3136 6276 3148
rect 6328 3136 6334 3188
rect 8205 3179 8263 3185
rect 8205 3145 8217 3179
rect 8251 3145 8263 3179
rect 8205 3139 8263 3145
rect 5169 3111 5227 3117
rect 5169 3077 5181 3111
rect 5215 3108 5227 3111
rect 7558 3108 7564 3120
rect 5215 3080 6132 3108
rect 7406 3080 7564 3108
rect 5215 3077 5227 3080
rect 5169 3071 5227 3077
rect 6104 3052 6132 3080
rect 7558 3068 7564 3080
rect 7616 3068 7622 3120
rect 7837 3111 7895 3117
rect 7837 3077 7849 3111
rect 7883 3108 7895 3111
rect 8220 3108 8248 3139
rect 9030 3136 9036 3188
rect 9088 3136 9094 3188
rect 11146 3136 11152 3188
rect 11204 3176 11210 3188
rect 11517 3179 11575 3185
rect 11517 3176 11529 3179
rect 11204 3148 11529 3176
rect 11204 3136 11210 3148
rect 11517 3145 11529 3148
rect 11563 3145 11575 3179
rect 13354 3176 13360 3188
rect 11517 3139 11575 3145
rect 12406 3148 13360 3176
rect 7883 3080 8248 3108
rect 7883 3077 7895 3080
rect 7837 3071 7895 3077
rect 4706 3000 4712 3052
rect 4764 3000 4770 3052
rect 4801 3043 4859 3049
rect 4801 3009 4813 3043
rect 4847 3040 4859 3043
rect 5445 3043 5503 3049
rect 5445 3040 5457 3043
rect 4847 3012 5457 3040
rect 4847 3009 4859 3012
rect 4801 3003 4859 3009
rect 5445 3009 5457 3012
rect 5491 3009 5503 3043
rect 5445 3003 5503 3009
rect 5350 2932 5356 2984
rect 5408 2932 5414 2984
rect 5460 2972 5488 3003
rect 5718 3000 5724 3052
rect 5776 3040 5782 3052
rect 5905 3043 5963 3049
rect 5905 3040 5917 3043
rect 5776 3012 5917 3040
rect 5776 3000 5782 3012
rect 5905 3009 5917 3012
rect 5951 3009 5963 3043
rect 5905 3003 5963 3009
rect 6086 3000 6092 3052
rect 6144 3000 6150 3052
rect 8113 3043 8171 3049
rect 8113 3009 8125 3043
rect 8159 3040 8171 3043
rect 8202 3040 8208 3052
rect 8159 3012 8208 3040
rect 8159 3009 8171 3012
rect 8113 3003 8171 3009
rect 8202 3000 8208 3012
rect 8260 3000 8266 3052
rect 8573 3043 8631 3049
rect 8573 3009 8585 3043
rect 8619 3040 8631 3043
rect 9048 3040 9076 3136
rect 11606 3108 11612 3120
rect 10074 3080 11612 3108
rect 11606 3068 11612 3080
rect 11664 3068 11670 3120
rect 12161 3111 12219 3117
rect 12161 3077 12173 3111
rect 12207 3108 12219 3111
rect 12406 3108 12434 3148
rect 13354 3136 13360 3148
rect 13412 3136 13418 3188
rect 14642 3136 14648 3188
rect 14700 3136 14706 3188
rect 15289 3179 15347 3185
rect 15289 3145 15301 3179
rect 15335 3176 15347 3179
rect 16574 3176 16580 3188
rect 15335 3148 16580 3176
rect 15335 3145 15347 3148
rect 15289 3139 15347 3145
rect 16574 3136 16580 3148
rect 16632 3136 16638 3188
rect 12207 3080 12480 3108
rect 12207 3077 12219 3080
rect 12161 3071 12219 3077
rect 8619 3012 9076 3040
rect 10781 3043 10839 3049
rect 8619 3009 8631 3012
rect 8573 3003 8631 3009
rect 10781 3009 10793 3043
rect 10827 3040 10839 3043
rect 11514 3040 11520 3052
rect 10827 3012 11520 3040
rect 10827 3009 10839 3012
rect 10781 3003 10839 3009
rect 11514 3000 11520 3012
rect 11572 3000 11578 3052
rect 11701 3043 11759 3049
rect 11701 3009 11713 3043
rect 11747 3040 11759 3043
rect 12250 3040 12256 3052
rect 11747 3012 12256 3040
rect 11747 3009 11759 3012
rect 11701 3003 11759 3009
rect 12250 3000 12256 3012
rect 12308 3000 12314 3052
rect 12452 3049 12480 3080
rect 13630 3068 13636 3120
rect 13688 3068 13694 3120
rect 14090 3068 14096 3120
rect 14148 3068 14154 3120
rect 15746 3108 15752 3120
rect 14844 3080 15752 3108
rect 12437 3043 12495 3049
rect 12437 3009 12449 3043
rect 12483 3009 12495 3043
rect 12437 3003 12495 3009
rect 14369 3043 14427 3049
rect 14369 3009 14381 3043
rect 14415 3040 14427 3043
rect 14458 3040 14464 3052
rect 14415 3012 14464 3040
rect 14415 3009 14427 3012
rect 14369 3003 14427 3009
rect 14458 3000 14464 3012
rect 14516 3000 14522 3052
rect 14844 3049 14872 3080
rect 15746 3068 15752 3080
rect 15804 3068 15810 3120
rect 14829 3043 14887 3049
rect 14829 3009 14841 3043
rect 14875 3009 14887 3043
rect 14829 3003 14887 3009
rect 14921 3043 14979 3049
rect 14921 3009 14933 3043
rect 14967 3040 14979 3043
rect 15194 3040 15200 3052
rect 14967 3012 15200 3040
rect 14967 3009 14979 3012
rect 14921 3003 14979 3009
rect 15194 3000 15200 3012
rect 15252 3000 15258 3052
rect 15654 3000 15660 3052
rect 15712 3000 15718 3052
rect 17034 3000 17040 3052
rect 17092 3000 17098 3052
rect 6365 2975 6423 2981
rect 6365 2972 6377 2975
rect 5460 2944 6377 2972
rect 6365 2941 6377 2944
rect 6411 2941 6423 2975
rect 6365 2935 6423 2941
rect 8662 2932 8668 2984
rect 8720 2932 8726 2984
rect 10505 2975 10563 2981
rect 10505 2941 10517 2975
rect 10551 2972 10563 2975
rect 11793 2975 11851 2981
rect 10551 2944 10732 2972
rect 10551 2941 10563 2944
rect 10505 2935 10563 2941
rect 10704 2904 10732 2944
rect 11793 2941 11805 2975
rect 11839 2972 11851 2975
rect 11882 2972 11888 2984
rect 11839 2944 11888 2972
rect 11839 2941 11851 2944
rect 11793 2935 11851 2941
rect 11882 2932 11888 2944
rect 11940 2972 11946 2984
rect 11940 2944 12434 2972
rect 11940 2932 11946 2944
rect 11514 2904 11520 2916
rect 10704 2876 11520 2904
rect 11514 2864 11520 2876
rect 11572 2864 11578 2916
rect 12406 2904 12434 2944
rect 12621 2907 12679 2913
rect 12621 2904 12633 2907
rect 12406 2876 12633 2904
rect 12621 2873 12633 2876
rect 12667 2873 12679 2907
rect 12621 2867 12679 2873
rect 15378 2864 15384 2916
rect 15436 2904 15442 2916
rect 15473 2907 15531 2913
rect 15473 2904 15485 2907
rect 15436 2876 15485 2904
rect 15436 2864 15442 2876
rect 15473 2873 15485 2876
rect 15519 2873 15531 2907
rect 15473 2867 15531 2873
rect 15562 2864 15568 2916
rect 15620 2904 15626 2916
rect 16853 2907 16911 2913
rect 16853 2904 16865 2907
rect 15620 2876 16865 2904
rect 15620 2864 15626 2876
rect 16853 2873 16865 2876
rect 16899 2873 16911 2907
rect 16853 2867 16911 2873
rect 5350 2796 5356 2848
rect 5408 2836 5414 2848
rect 5997 2839 6055 2845
rect 5997 2836 6009 2839
rect 5408 2808 6009 2836
rect 5408 2796 5414 2808
rect 5997 2805 6009 2808
rect 6043 2805 6055 2839
rect 5997 2799 6055 2805
rect 11974 2796 11980 2848
rect 12032 2836 12038 2848
rect 12345 2839 12403 2845
rect 12345 2836 12357 2839
rect 12032 2808 12357 2836
rect 12032 2796 12038 2808
rect 12345 2805 12357 2808
rect 12391 2805 12403 2839
rect 12345 2799 12403 2805
rect 1104 2746 17388 2768
rect 1104 2694 2985 2746
rect 3037 2694 3049 2746
rect 3101 2694 3113 2746
rect 3165 2694 3177 2746
rect 3229 2694 3241 2746
rect 3293 2694 7056 2746
rect 7108 2694 7120 2746
rect 7172 2694 7184 2746
rect 7236 2694 7248 2746
rect 7300 2694 7312 2746
rect 7364 2694 11127 2746
rect 11179 2694 11191 2746
rect 11243 2694 11255 2746
rect 11307 2694 11319 2746
rect 11371 2694 11383 2746
rect 11435 2694 15198 2746
rect 15250 2694 15262 2746
rect 15314 2694 15326 2746
rect 15378 2694 15390 2746
rect 15442 2694 15454 2746
rect 15506 2694 17388 2746
rect 1104 2672 17388 2694
rect 5442 2592 5448 2644
rect 5500 2592 5506 2644
rect 6822 2592 6828 2644
rect 6880 2632 6886 2644
rect 7377 2635 7435 2641
rect 7377 2632 7389 2635
rect 6880 2604 7389 2632
rect 6880 2592 6886 2604
rect 7377 2601 7389 2604
rect 7423 2601 7435 2635
rect 7377 2595 7435 2601
rect 8294 2592 8300 2644
rect 8352 2632 8358 2644
rect 8481 2635 8539 2641
rect 8481 2632 8493 2635
rect 8352 2604 8493 2632
rect 8352 2592 8358 2604
rect 8481 2601 8493 2604
rect 8527 2601 8539 2635
rect 8481 2595 8539 2601
rect 9953 2635 10011 2641
rect 9953 2601 9965 2635
rect 9999 2632 10011 2635
rect 10134 2632 10140 2644
rect 9999 2604 10140 2632
rect 9999 2601 10011 2604
rect 9953 2595 10011 2601
rect 10134 2592 10140 2604
rect 10192 2592 10198 2644
rect 10226 2592 10232 2644
rect 10284 2632 10290 2644
rect 10597 2635 10655 2641
rect 10597 2632 10609 2635
rect 10284 2604 10609 2632
rect 10284 2592 10290 2604
rect 10597 2601 10609 2604
rect 10643 2601 10655 2635
rect 10597 2595 10655 2601
rect 11241 2635 11299 2641
rect 11241 2601 11253 2635
rect 11287 2632 11299 2635
rect 11606 2632 11612 2644
rect 11287 2604 11612 2632
rect 11287 2601 11299 2604
rect 11241 2595 11299 2601
rect 11606 2592 11612 2604
rect 11664 2592 11670 2644
rect 13173 2635 13231 2641
rect 13173 2601 13185 2635
rect 13219 2632 13231 2635
rect 13446 2632 13452 2644
rect 13219 2604 13452 2632
rect 13219 2601 13231 2604
rect 13173 2595 13231 2601
rect 13446 2592 13452 2604
rect 13504 2592 13510 2644
rect 11514 2524 11520 2576
rect 11572 2524 11578 2576
rect 11974 2456 11980 2508
rect 12032 2456 12038 2508
rect 5166 2388 5172 2440
rect 5224 2428 5230 2440
rect 5261 2431 5319 2437
rect 5261 2428 5273 2431
rect 5224 2400 5273 2428
rect 5224 2388 5230 2400
rect 5261 2397 5273 2400
rect 5307 2397 5319 2431
rect 5261 2391 5319 2397
rect 7098 2388 7104 2440
rect 7156 2428 7162 2440
rect 7193 2431 7251 2437
rect 7193 2428 7205 2431
rect 7156 2400 7205 2428
rect 7156 2388 7162 2400
rect 7193 2397 7205 2400
rect 7239 2397 7251 2431
rect 7193 2391 7251 2397
rect 8386 2388 8392 2440
rect 8444 2428 8450 2440
rect 8665 2431 8723 2437
rect 8665 2428 8677 2431
rect 8444 2400 8677 2428
rect 8444 2388 8450 2400
rect 8665 2397 8677 2400
rect 8711 2397 8723 2431
rect 8665 2391 8723 2397
rect 9674 2388 9680 2440
rect 9732 2428 9738 2440
rect 9769 2431 9827 2437
rect 9769 2428 9781 2431
rect 9732 2400 9781 2428
rect 9732 2388 9738 2400
rect 9769 2397 9781 2400
rect 9815 2397 9827 2431
rect 9769 2391 9827 2397
rect 10318 2388 10324 2440
rect 10376 2428 10382 2440
rect 10413 2431 10471 2437
rect 10413 2428 10425 2431
rect 10376 2400 10425 2428
rect 10376 2388 10382 2400
rect 10413 2397 10425 2400
rect 10459 2397 10471 2431
rect 10413 2391 10471 2397
rect 10962 2388 10968 2440
rect 11020 2428 11026 2440
rect 11057 2431 11115 2437
rect 11057 2428 11069 2431
rect 11020 2400 11069 2428
rect 11020 2388 11026 2400
rect 11057 2397 11069 2400
rect 11103 2397 11115 2431
rect 11057 2391 11115 2397
rect 11882 2388 11888 2440
rect 11940 2388 11946 2440
rect 12894 2388 12900 2440
rect 12952 2428 12958 2440
rect 12989 2431 13047 2437
rect 12989 2428 13001 2431
rect 12952 2400 13001 2428
rect 12952 2388 12958 2400
rect 12989 2397 13001 2400
rect 13035 2397 13047 2431
rect 12989 2391 13047 2397
rect 1104 2202 17388 2224
rect 1104 2150 3645 2202
rect 3697 2150 3709 2202
rect 3761 2150 3773 2202
rect 3825 2150 3837 2202
rect 3889 2150 3901 2202
rect 3953 2150 7716 2202
rect 7768 2150 7780 2202
rect 7832 2150 7844 2202
rect 7896 2150 7908 2202
rect 7960 2150 7972 2202
rect 8024 2150 11787 2202
rect 11839 2150 11851 2202
rect 11903 2150 11915 2202
rect 11967 2150 11979 2202
rect 12031 2150 12043 2202
rect 12095 2150 15858 2202
rect 15910 2150 15922 2202
rect 15974 2150 15986 2202
rect 16038 2150 16050 2202
rect 16102 2150 16114 2202
rect 16166 2150 17388 2202
rect 1104 2128 17388 2150
<< via1 >>
rect 2985 17926 3037 17978
rect 3049 17926 3101 17978
rect 3113 17926 3165 17978
rect 3177 17926 3229 17978
rect 3241 17926 3293 17978
rect 7056 17926 7108 17978
rect 7120 17926 7172 17978
rect 7184 17926 7236 17978
rect 7248 17926 7300 17978
rect 7312 17926 7364 17978
rect 11127 17926 11179 17978
rect 11191 17926 11243 17978
rect 11255 17926 11307 17978
rect 11319 17926 11371 17978
rect 11383 17926 11435 17978
rect 15198 17926 15250 17978
rect 15262 17926 15314 17978
rect 15326 17926 15378 17978
rect 15390 17926 15442 17978
rect 15454 17926 15506 17978
rect 9588 17824 9640 17876
rect 12348 17824 12400 17876
rect 5080 17756 5132 17808
rect 8944 17756 8996 17808
rect 5172 17688 5224 17740
rect 4068 17620 4120 17672
rect 5448 17620 5500 17672
rect 5080 17595 5132 17604
rect 5080 17561 5089 17595
rect 5089 17561 5123 17595
rect 5123 17561 5132 17595
rect 5080 17552 5132 17561
rect 5264 17595 5316 17604
rect 5264 17561 5273 17595
rect 5273 17561 5307 17595
rect 5307 17561 5316 17595
rect 5264 17552 5316 17561
rect 8392 17620 8444 17672
rect 9036 17688 9088 17740
rect 9404 17688 9456 17740
rect 8944 17663 8996 17672
rect 8944 17629 8953 17663
rect 8953 17629 8987 17663
rect 8987 17629 8996 17663
rect 8944 17620 8996 17629
rect 9128 17620 9180 17672
rect 5908 17552 5960 17604
rect 9772 17620 9824 17672
rect 10968 17620 11020 17672
rect 12256 17620 12308 17672
rect 10048 17595 10100 17604
rect 10048 17561 10057 17595
rect 10057 17561 10091 17595
rect 10091 17561 10100 17595
rect 10048 17552 10100 17561
rect 13084 17552 13136 17604
rect 5540 17484 5592 17536
rect 8484 17527 8536 17536
rect 8484 17493 8493 17527
rect 8493 17493 8527 17527
rect 8527 17493 8536 17527
rect 8484 17484 8536 17493
rect 8576 17527 8628 17536
rect 8576 17493 8585 17527
rect 8585 17493 8619 17527
rect 8619 17493 8628 17527
rect 8576 17484 8628 17493
rect 8668 17484 8720 17536
rect 9220 17484 9272 17536
rect 9404 17527 9456 17536
rect 9404 17493 9413 17527
rect 9413 17493 9447 17527
rect 9447 17493 9456 17527
rect 9404 17484 9456 17493
rect 9496 17484 9548 17536
rect 11520 17484 11572 17536
rect 12532 17527 12584 17536
rect 12532 17493 12541 17527
rect 12541 17493 12575 17527
rect 12575 17493 12584 17527
rect 12532 17484 12584 17493
rect 3645 17382 3697 17434
rect 3709 17382 3761 17434
rect 3773 17382 3825 17434
rect 3837 17382 3889 17434
rect 3901 17382 3953 17434
rect 7716 17382 7768 17434
rect 7780 17382 7832 17434
rect 7844 17382 7896 17434
rect 7908 17382 7960 17434
rect 7972 17382 8024 17434
rect 11787 17382 11839 17434
rect 11851 17382 11903 17434
rect 11915 17382 11967 17434
rect 11979 17382 12031 17434
rect 12043 17382 12095 17434
rect 15858 17382 15910 17434
rect 15922 17382 15974 17434
rect 15986 17382 16038 17434
rect 16050 17382 16102 17434
rect 16114 17382 16166 17434
rect 5908 17323 5960 17332
rect 5908 17289 5917 17323
rect 5917 17289 5951 17323
rect 5951 17289 5960 17323
rect 5908 17280 5960 17289
rect 8944 17280 8996 17332
rect 9128 17280 9180 17332
rect 4160 17212 4212 17264
rect 5540 17212 5592 17264
rect 9312 17280 9364 17332
rect 848 17144 900 17196
rect 5448 17187 5500 17196
rect 5448 17153 5457 17187
rect 5457 17153 5491 17187
rect 5491 17153 5500 17187
rect 5448 17144 5500 17153
rect 6000 17144 6052 17196
rect 3424 17119 3476 17128
rect 3424 17085 3433 17119
rect 3433 17085 3467 17119
rect 3467 17085 3476 17119
rect 3424 17076 3476 17085
rect 6276 17076 6328 17128
rect 6552 17076 6604 17128
rect 6736 17187 6788 17196
rect 6736 17153 6745 17187
rect 6745 17153 6779 17187
rect 6779 17153 6788 17187
rect 6736 17144 6788 17153
rect 8392 17144 8444 17196
rect 9404 17144 9456 17196
rect 9588 17187 9640 17196
rect 9588 17153 9597 17187
rect 9597 17153 9631 17187
rect 9631 17153 9640 17187
rect 9588 17144 9640 17153
rect 9220 17076 9272 17128
rect 9864 17119 9916 17128
rect 9864 17085 9873 17119
rect 9873 17085 9907 17119
rect 9907 17085 9916 17119
rect 9864 17076 9916 17085
rect 10876 17076 10928 17128
rect 12992 17119 13044 17128
rect 12992 17085 13001 17119
rect 13001 17085 13035 17119
rect 13035 17085 13044 17119
rect 12992 17076 13044 17085
rect 1584 16983 1636 16992
rect 1584 16949 1593 16983
rect 1593 16949 1627 16983
rect 1627 16949 1636 16983
rect 1584 16940 1636 16949
rect 5264 16940 5316 16992
rect 6092 16940 6144 16992
rect 6460 16983 6512 16992
rect 6460 16949 6469 16983
rect 6469 16949 6503 16983
rect 6503 16949 6512 16983
rect 6460 16940 6512 16949
rect 9128 16940 9180 16992
rect 9588 16940 9640 16992
rect 10324 16940 10376 16992
rect 12348 16940 12400 16992
rect 2985 16838 3037 16890
rect 3049 16838 3101 16890
rect 3113 16838 3165 16890
rect 3177 16838 3229 16890
rect 3241 16838 3293 16890
rect 7056 16838 7108 16890
rect 7120 16838 7172 16890
rect 7184 16838 7236 16890
rect 7248 16838 7300 16890
rect 7312 16838 7364 16890
rect 11127 16838 11179 16890
rect 11191 16838 11243 16890
rect 11255 16838 11307 16890
rect 11319 16838 11371 16890
rect 11383 16838 11435 16890
rect 15198 16838 15250 16890
rect 15262 16838 15314 16890
rect 15326 16838 15378 16890
rect 15390 16838 15442 16890
rect 15454 16838 15506 16890
rect 5448 16736 5500 16788
rect 6000 16736 6052 16788
rect 9220 16779 9272 16788
rect 9220 16745 9229 16779
rect 9229 16745 9263 16779
rect 9263 16745 9272 16779
rect 9220 16736 9272 16745
rect 9864 16779 9916 16788
rect 9864 16745 9873 16779
rect 9873 16745 9907 16779
rect 9907 16745 9916 16779
rect 9864 16736 9916 16745
rect 12992 16736 13044 16788
rect 10048 16668 10100 16720
rect 6092 16600 6144 16652
rect 6460 16643 6512 16652
rect 6460 16609 6469 16643
rect 6469 16609 6503 16643
rect 6503 16609 6512 16643
rect 6460 16600 6512 16609
rect 9496 16643 9548 16652
rect 9496 16609 9505 16643
rect 9505 16609 9539 16643
rect 9539 16609 9548 16643
rect 9496 16600 9548 16609
rect 11704 16600 11756 16652
rect 1584 16575 1636 16584
rect 1584 16541 1593 16575
rect 1593 16541 1627 16575
rect 1627 16541 1636 16575
rect 1584 16532 1636 16541
rect 5080 16575 5132 16584
rect 5080 16541 5089 16575
rect 5089 16541 5123 16575
rect 5123 16541 5132 16575
rect 5080 16532 5132 16541
rect 5264 16532 5316 16584
rect 8392 16532 8444 16584
rect 8944 16575 8996 16584
rect 8944 16541 8953 16575
rect 8953 16541 8987 16575
rect 8987 16541 8996 16575
rect 8944 16532 8996 16541
rect 9036 16532 9088 16584
rect 1584 16396 1636 16448
rect 6000 16464 6052 16516
rect 8208 16464 8260 16516
rect 9312 16532 9364 16584
rect 11612 16532 11664 16584
rect 5080 16396 5132 16448
rect 8116 16396 8168 16448
rect 3645 16294 3697 16346
rect 3709 16294 3761 16346
rect 3773 16294 3825 16346
rect 3837 16294 3889 16346
rect 3901 16294 3953 16346
rect 7716 16294 7768 16346
rect 7780 16294 7832 16346
rect 7844 16294 7896 16346
rect 7908 16294 7960 16346
rect 7972 16294 8024 16346
rect 11787 16294 11839 16346
rect 11851 16294 11903 16346
rect 11915 16294 11967 16346
rect 11979 16294 12031 16346
rect 12043 16294 12095 16346
rect 15858 16294 15910 16346
rect 15922 16294 15974 16346
rect 15986 16294 16038 16346
rect 16050 16294 16102 16346
rect 16114 16294 16166 16346
rect 4160 16124 4212 16176
rect 5172 16124 5224 16176
rect 3332 16099 3384 16108
rect 3332 16065 3341 16099
rect 3341 16065 3375 16099
rect 3375 16065 3384 16099
rect 3332 16056 3384 16065
rect 3516 16099 3568 16108
rect 3516 16065 3525 16099
rect 3525 16065 3559 16099
rect 3559 16065 3568 16099
rect 3516 16056 3568 16065
rect 1400 16031 1452 16040
rect 1400 15997 1409 16031
rect 1409 15997 1443 16031
rect 1443 15997 1452 16031
rect 1400 15988 1452 15997
rect 1676 16031 1728 16040
rect 1676 15997 1685 16031
rect 1685 15997 1719 16031
rect 1719 15997 1728 16031
rect 1676 15988 1728 15997
rect 2780 15852 2832 15904
rect 3884 15852 3936 15904
rect 2985 15750 3037 15802
rect 3049 15750 3101 15802
rect 3113 15750 3165 15802
rect 3177 15750 3229 15802
rect 3241 15750 3293 15802
rect 7056 15750 7108 15802
rect 7120 15750 7172 15802
rect 7184 15750 7236 15802
rect 7248 15750 7300 15802
rect 7312 15750 7364 15802
rect 11127 15750 11179 15802
rect 11191 15750 11243 15802
rect 11255 15750 11307 15802
rect 11319 15750 11371 15802
rect 11383 15750 11435 15802
rect 15198 15750 15250 15802
rect 15262 15750 15314 15802
rect 15326 15750 15378 15802
rect 15390 15750 15442 15802
rect 15454 15750 15506 15802
rect 1676 15648 1728 15700
rect 3240 15648 3292 15700
rect 4068 15648 4120 15700
rect 1400 15580 1452 15632
rect 3424 15580 3476 15632
rect 6276 15648 6328 15700
rect 11704 15691 11756 15700
rect 11704 15657 11713 15691
rect 11713 15657 11747 15691
rect 11747 15657 11756 15691
rect 11704 15648 11756 15657
rect 1032 15444 1084 15496
rect 3240 15512 3292 15564
rect 3884 15555 3936 15564
rect 3884 15521 3893 15555
rect 3893 15521 3927 15555
rect 3927 15521 3936 15555
rect 3884 15512 3936 15521
rect 5264 15512 5316 15564
rect 8208 15512 8260 15564
rect 1584 15419 1636 15428
rect 1584 15385 1593 15419
rect 1593 15385 1627 15419
rect 1627 15385 1636 15419
rect 1584 15376 1636 15385
rect 2872 15444 2924 15496
rect 2964 15487 3016 15496
rect 2964 15453 2973 15487
rect 2973 15453 3007 15487
rect 3007 15453 3016 15487
rect 2964 15444 3016 15453
rect 3976 15487 4028 15496
rect 3976 15453 3985 15487
rect 3985 15453 4019 15487
rect 4019 15453 4028 15487
rect 3976 15444 4028 15453
rect 7564 15444 7616 15496
rect 2688 15419 2740 15428
rect 2688 15385 2697 15419
rect 2697 15385 2731 15419
rect 2731 15385 2740 15419
rect 2688 15376 2740 15385
rect 3332 15308 3384 15360
rect 5172 15376 5224 15428
rect 7472 15376 7524 15428
rect 8484 15487 8536 15496
rect 8484 15453 8493 15487
rect 8493 15453 8527 15487
rect 8527 15453 8536 15487
rect 8484 15444 8536 15453
rect 9312 15487 9364 15496
rect 9312 15453 9321 15487
rect 9321 15453 9355 15487
rect 9355 15453 9364 15487
rect 9312 15444 9364 15453
rect 8300 15419 8352 15428
rect 8300 15385 8309 15419
rect 8309 15385 8343 15419
rect 8343 15385 8352 15419
rect 8300 15376 8352 15385
rect 9588 15419 9640 15428
rect 9588 15385 9597 15419
rect 9597 15385 9631 15419
rect 9631 15385 9640 15419
rect 9588 15376 9640 15385
rect 10876 15376 10928 15428
rect 11704 15444 11756 15496
rect 12624 15580 12676 15632
rect 12532 15444 12584 15496
rect 13084 15487 13136 15496
rect 13084 15453 13093 15487
rect 13093 15453 13127 15487
rect 13127 15453 13136 15487
rect 13084 15444 13136 15453
rect 7012 15308 7064 15360
rect 9404 15308 9456 15360
rect 11612 15308 11664 15360
rect 12256 15419 12308 15428
rect 12256 15385 12265 15419
rect 12265 15385 12299 15419
rect 12299 15385 12308 15419
rect 12256 15376 12308 15385
rect 14924 15512 14976 15564
rect 16580 15444 16632 15496
rect 17040 15487 17092 15496
rect 17040 15453 17049 15487
rect 17049 15453 17083 15487
rect 17083 15453 17092 15487
rect 17040 15444 17092 15453
rect 14924 15419 14976 15428
rect 14924 15385 14933 15419
rect 14933 15385 14967 15419
rect 14967 15385 14976 15419
rect 14924 15376 14976 15385
rect 12164 15308 12216 15360
rect 13268 15351 13320 15360
rect 13268 15317 13277 15351
rect 13277 15317 13311 15351
rect 13311 15317 13320 15351
rect 13268 15308 13320 15317
rect 14188 15351 14240 15360
rect 14188 15317 14197 15351
rect 14197 15317 14231 15351
rect 14231 15317 14240 15351
rect 14188 15308 14240 15317
rect 14556 15351 14608 15360
rect 14556 15317 14565 15351
rect 14565 15317 14599 15351
rect 14599 15317 14608 15351
rect 14556 15308 14608 15317
rect 14740 15351 14792 15360
rect 14740 15317 14749 15351
rect 14749 15317 14783 15351
rect 14783 15317 14792 15351
rect 14740 15308 14792 15317
rect 16856 15351 16908 15360
rect 16856 15317 16865 15351
rect 16865 15317 16899 15351
rect 16899 15317 16908 15351
rect 16856 15308 16908 15317
rect 3645 15206 3697 15258
rect 3709 15206 3761 15258
rect 3773 15206 3825 15258
rect 3837 15206 3889 15258
rect 3901 15206 3953 15258
rect 7716 15206 7768 15258
rect 7780 15206 7832 15258
rect 7844 15206 7896 15258
rect 7908 15206 7960 15258
rect 7972 15206 8024 15258
rect 11787 15206 11839 15258
rect 11851 15206 11903 15258
rect 11915 15206 11967 15258
rect 11979 15206 12031 15258
rect 12043 15206 12095 15258
rect 15858 15206 15910 15258
rect 15922 15206 15974 15258
rect 15986 15206 16038 15258
rect 16050 15206 16102 15258
rect 16114 15206 16166 15258
rect 2964 15104 3016 15156
rect 3516 15147 3568 15156
rect 3516 15113 3525 15147
rect 3525 15113 3559 15147
rect 3559 15113 3568 15147
rect 3516 15104 3568 15113
rect 8300 15104 8352 15156
rect 9588 15104 9640 15156
rect 14924 15104 14976 15156
rect 2780 15036 2832 15088
rect 2872 14968 2924 15020
rect 7012 15079 7064 15088
rect 7012 15045 7021 15079
rect 7021 15045 7055 15079
rect 7055 15045 7064 15079
rect 7012 15036 7064 15045
rect 8392 15036 8444 15088
rect 6092 14968 6144 15020
rect 3516 14900 3568 14952
rect 5080 14900 5132 14952
rect 7472 14900 7524 14952
rect 15660 15036 15712 15088
rect 7380 14764 7432 14816
rect 7564 14764 7616 14816
rect 9404 15011 9456 15020
rect 9404 14977 9413 15011
rect 9413 14977 9447 15011
rect 9447 14977 9456 15011
rect 9404 14968 9456 14977
rect 12900 14968 12952 15020
rect 13268 14968 13320 15020
rect 11888 14900 11940 14952
rect 14096 14900 14148 14952
rect 14372 14900 14424 14952
rect 14924 14900 14976 14952
rect 11796 14764 11848 14816
rect 12256 14764 12308 14816
rect 15568 14764 15620 14816
rect 2985 14662 3037 14714
rect 3049 14662 3101 14714
rect 3113 14662 3165 14714
rect 3177 14662 3229 14714
rect 3241 14662 3293 14714
rect 7056 14662 7108 14714
rect 7120 14662 7172 14714
rect 7184 14662 7236 14714
rect 7248 14662 7300 14714
rect 7312 14662 7364 14714
rect 11127 14662 11179 14714
rect 11191 14662 11243 14714
rect 11255 14662 11307 14714
rect 11319 14662 11371 14714
rect 11383 14662 11435 14714
rect 15198 14662 15250 14714
rect 15262 14662 15314 14714
rect 15326 14662 15378 14714
rect 15390 14662 15442 14714
rect 15454 14662 15506 14714
rect 3976 14560 4028 14612
rect 7472 14560 7524 14612
rect 11888 14603 11940 14612
rect 11888 14569 11897 14603
rect 11897 14569 11931 14603
rect 11931 14569 11940 14603
rect 11888 14560 11940 14569
rect 14096 14603 14148 14612
rect 14096 14569 14105 14603
rect 14105 14569 14139 14603
rect 14139 14569 14148 14603
rect 14096 14560 14148 14569
rect 14924 14603 14976 14612
rect 14924 14569 14933 14603
rect 14933 14569 14967 14603
rect 14967 14569 14976 14603
rect 14924 14560 14976 14569
rect 17040 14603 17092 14612
rect 17040 14569 17049 14603
rect 17049 14569 17083 14603
rect 17083 14569 17092 14603
rect 17040 14560 17092 14569
rect 7380 14492 7432 14544
rect 8668 14492 8720 14544
rect 11796 14492 11848 14544
rect 12348 14492 12400 14544
rect 5264 14424 5316 14476
rect 6092 14424 6144 14476
rect 7564 14424 7616 14476
rect 10232 14467 10284 14476
rect 10232 14433 10241 14467
rect 10241 14433 10275 14467
rect 10275 14433 10284 14467
rect 10232 14424 10284 14433
rect 11612 14467 11664 14476
rect 11612 14433 11621 14467
rect 11621 14433 11655 14467
rect 11655 14433 11664 14467
rect 11612 14424 11664 14433
rect 11704 14467 11756 14476
rect 11704 14433 11713 14467
rect 11713 14433 11747 14467
rect 11747 14433 11756 14467
rect 11704 14424 11756 14433
rect 14556 14424 14608 14476
rect 14740 14467 14792 14476
rect 14740 14433 14749 14467
rect 14749 14433 14783 14467
rect 14783 14433 14792 14467
rect 14740 14424 14792 14433
rect 5172 14288 5224 14340
rect 6092 14331 6144 14340
rect 6092 14297 6101 14331
rect 6101 14297 6135 14331
rect 6135 14297 6144 14331
rect 6092 14288 6144 14297
rect 7564 14288 7616 14340
rect 8300 14356 8352 14408
rect 8484 14356 8536 14408
rect 10324 14356 10376 14408
rect 12164 14356 12216 14408
rect 12256 14399 12308 14408
rect 12256 14365 12265 14399
rect 12265 14365 12299 14399
rect 12299 14365 12308 14399
rect 12256 14356 12308 14365
rect 12532 14399 12584 14408
rect 12532 14365 12541 14399
rect 12541 14365 12575 14399
rect 12575 14365 12584 14399
rect 12532 14356 12584 14365
rect 13268 14356 13320 14408
rect 14372 14399 14424 14408
rect 14372 14365 14381 14399
rect 14381 14365 14415 14399
rect 14415 14365 14424 14399
rect 14372 14356 14424 14365
rect 15568 14467 15620 14476
rect 15568 14433 15577 14467
rect 15577 14433 15611 14467
rect 15611 14433 15620 14467
rect 15568 14424 15620 14433
rect 8668 14220 8720 14272
rect 12440 14331 12492 14340
rect 12440 14297 12449 14331
rect 12449 14297 12483 14331
rect 12483 14297 12492 14331
rect 12440 14288 12492 14297
rect 14188 14288 14240 14340
rect 14280 14288 14332 14340
rect 15660 14288 15712 14340
rect 3645 14118 3697 14170
rect 3709 14118 3761 14170
rect 3773 14118 3825 14170
rect 3837 14118 3889 14170
rect 3901 14118 3953 14170
rect 7716 14118 7768 14170
rect 7780 14118 7832 14170
rect 7844 14118 7896 14170
rect 7908 14118 7960 14170
rect 7972 14118 8024 14170
rect 11787 14118 11839 14170
rect 11851 14118 11903 14170
rect 11915 14118 11967 14170
rect 11979 14118 12031 14170
rect 12043 14118 12095 14170
rect 15858 14118 15910 14170
rect 15922 14118 15974 14170
rect 15986 14118 16038 14170
rect 16050 14118 16102 14170
rect 16114 14118 16166 14170
rect 2780 14016 2832 14068
rect 6092 14016 6144 14068
rect 7564 14016 7616 14068
rect 8392 14016 8444 14068
rect 10232 14059 10284 14068
rect 10232 14025 10241 14059
rect 10241 14025 10275 14059
rect 10275 14025 10284 14059
rect 10232 14016 10284 14025
rect 14372 14016 14424 14068
rect 16580 14016 16632 14068
rect 15660 13948 15712 14000
rect 1400 13923 1452 13932
rect 1400 13889 1409 13923
rect 1409 13889 1443 13923
rect 1443 13889 1452 13923
rect 1400 13880 1452 13889
rect 5540 13880 5592 13932
rect 10140 13880 10192 13932
rect 10416 13923 10468 13932
rect 10416 13889 10425 13923
rect 10425 13889 10459 13923
rect 10459 13889 10468 13923
rect 10416 13880 10468 13889
rect 17040 13923 17092 13932
rect 17040 13889 17049 13923
rect 17049 13889 17083 13923
rect 17083 13889 17092 13923
rect 17040 13880 17092 13889
rect 5356 13855 5408 13864
rect 5356 13821 5365 13855
rect 5365 13821 5399 13855
rect 5399 13821 5408 13855
rect 5356 13812 5408 13821
rect 14280 13812 14332 13864
rect 16212 13719 16264 13728
rect 16212 13685 16233 13719
rect 16233 13685 16264 13719
rect 16212 13676 16264 13685
rect 2985 13574 3037 13626
rect 3049 13574 3101 13626
rect 3113 13574 3165 13626
rect 3177 13574 3229 13626
rect 3241 13574 3293 13626
rect 7056 13574 7108 13626
rect 7120 13574 7172 13626
rect 7184 13574 7236 13626
rect 7248 13574 7300 13626
rect 7312 13574 7364 13626
rect 11127 13574 11179 13626
rect 11191 13574 11243 13626
rect 11255 13574 11307 13626
rect 11319 13574 11371 13626
rect 11383 13574 11435 13626
rect 15198 13574 15250 13626
rect 15262 13574 15314 13626
rect 15326 13574 15378 13626
rect 15390 13574 15442 13626
rect 15454 13574 15506 13626
rect 5356 13472 5408 13524
rect 2780 13336 2832 13388
rect 848 13268 900 13320
rect 3332 13336 3384 13388
rect 3976 13268 4028 13320
rect 3240 13243 3292 13252
rect 3240 13209 3249 13243
rect 3249 13209 3283 13243
rect 3283 13209 3292 13243
rect 3240 13200 3292 13209
rect 2688 13175 2740 13184
rect 2688 13141 2697 13175
rect 2697 13141 2731 13175
rect 2731 13141 2740 13175
rect 2688 13132 2740 13141
rect 3424 13175 3476 13184
rect 3424 13141 3433 13175
rect 3433 13141 3467 13175
rect 3467 13141 3476 13175
rect 3424 13132 3476 13141
rect 3516 13132 3568 13184
rect 5540 13311 5592 13320
rect 5540 13277 5549 13311
rect 5549 13277 5583 13311
rect 5583 13277 5592 13311
rect 5540 13268 5592 13277
rect 6276 13311 6328 13320
rect 6276 13277 6285 13311
rect 6285 13277 6319 13311
rect 6319 13277 6328 13311
rect 6276 13268 6328 13277
rect 6368 13268 6420 13320
rect 6920 13311 6972 13320
rect 6920 13277 6929 13311
rect 6929 13277 6963 13311
rect 6963 13277 6972 13311
rect 6920 13268 6972 13277
rect 4712 13200 4764 13252
rect 7380 13268 7432 13320
rect 8116 13336 8168 13388
rect 10416 13404 10468 13456
rect 8576 13336 8628 13388
rect 10324 13336 10376 13388
rect 11612 13404 11664 13456
rect 12624 13404 12676 13456
rect 12440 13336 12492 13388
rect 8944 13200 8996 13252
rect 6368 13132 6420 13184
rect 6460 13175 6512 13184
rect 6460 13141 6469 13175
rect 6469 13141 6503 13175
rect 6503 13141 6512 13175
rect 6460 13132 6512 13141
rect 7564 13132 7616 13184
rect 9588 13132 9640 13184
rect 10140 13311 10192 13320
rect 10140 13277 10149 13311
rect 10149 13277 10183 13311
rect 10183 13277 10192 13311
rect 10140 13268 10192 13277
rect 11060 13311 11112 13320
rect 11060 13277 11069 13311
rect 11069 13277 11103 13311
rect 11103 13277 11112 13311
rect 11060 13268 11112 13277
rect 11428 13311 11480 13320
rect 11428 13277 11437 13311
rect 11437 13277 11471 13311
rect 11471 13277 11480 13311
rect 11428 13268 11480 13277
rect 10968 13200 11020 13252
rect 11612 13268 11664 13320
rect 13176 13311 13228 13320
rect 13176 13277 13185 13311
rect 13185 13277 13219 13311
rect 13219 13277 13228 13311
rect 13176 13268 13228 13277
rect 13544 13268 13596 13320
rect 17040 13311 17092 13320
rect 17040 13277 17049 13311
rect 17049 13277 17083 13311
rect 17083 13277 17092 13311
rect 17040 13268 17092 13277
rect 13728 13175 13780 13184
rect 13728 13141 13737 13175
rect 13737 13141 13771 13175
rect 13771 13141 13780 13175
rect 13728 13132 13780 13141
rect 3645 13030 3697 13082
rect 3709 13030 3761 13082
rect 3773 13030 3825 13082
rect 3837 13030 3889 13082
rect 3901 13030 3953 13082
rect 7716 13030 7768 13082
rect 7780 13030 7832 13082
rect 7844 13030 7896 13082
rect 7908 13030 7960 13082
rect 7972 13030 8024 13082
rect 11787 13030 11839 13082
rect 11851 13030 11903 13082
rect 11915 13030 11967 13082
rect 11979 13030 12031 13082
rect 12043 13030 12095 13082
rect 15858 13030 15910 13082
rect 15922 13030 15974 13082
rect 15986 13030 16038 13082
rect 16050 13030 16102 13082
rect 16114 13030 16166 13082
rect 3240 12928 3292 12980
rect 4712 12903 4764 12912
rect 4712 12869 4721 12903
rect 4721 12869 4755 12903
rect 4755 12869 4764 12903
rect 4712 12860 4764 12869
rect 6276 12928 6328 12980
rect 8944 12971 8996 12980
rect 8944 12937 8953 12971
rect 8953 12937 8987 12971
rect 8987 12937 8996 12971
rect 8944 12928 8996 12937
rect 10968 12928 11020 12980
rect 13176 12928 13228 12980
rect 13728 12928 13780 12980
rect 5172 12860 5224 12912
rect 8484 12860 8536 12912
rect 9588 12903 9640 12912
rect 9588 12869 9597 12903
rect 9597 12869 9631 12903
rect 9631 12869 9640 12903
rect 9588 12860 9640 12869
rect 10876 12860 10928 12912
rect 1400 12835 1452 12844
rect 1400 12801 1409 12835
rect 1409 12801 1443 12835
rect 1443 12801 1452 12835
rect 1400 12792 1452 12801
rect 2780 12792 2832 12844
rect 12900 12792 12952 12844
rect 13544 12835 13596 12844
rect 13544 12801 13553 12835
rect 13553 12801 13587 12835
rect 13587 12801 13596 12835
rect 13544 12792 13596 12801
rect 14280 12835 14332 12844
rect 14280 12801 14289 12835
rect 14289 12801 14323 12835
rect 14323 12801 14332 12835
rect 14280 12792 14332 12801
rect 15660 12792 15712 12844
rect 1676 12767 1728 12776
rect 1676 12733 1685 12767
rect 1685 12733 1719 12767
rect 1719 12733 1728 12767
rect 1676 12724 1728 12733
rect 2872 12724 2924 12776
rect 3332 12767 3384 12776
rect 3332 12733 3341 12767
rect 3341 12733 3375 12767
rect 3375 12733 3384 12767
rect 3332 12724 3384 12733
rect 4436 12767 4488 12776
rect 4436 12733 4445 12767
rect 4445 12733 4479 12767
rect 4479 12733 4488 12767
rect 4436 12724 4488 12733
rect 5264 12724 5316 12776
rect 6184 12724 6236 12776
rect 6828 12724 6880 12776
rect 7472 12767 7524 12776
rect 7472 12733 7481 12767
rect 7481 12733 7515 12767
rect 7515 12733 7524 12767
rect 7472 12724 7524 12733
rect 9312 12767 9364 12776
rect 9312 12733 9321 12767
rect 9321 12733 9355 12767
rect 9355 12733 9364 12767
rect 9312 12724 9364 12733
rect 11520 12767 11572 12776
rect 11520 12733 11529 12767
rect 11529 12733 11563 12767
rect 11563 12733 11572 12767
rect 11520 12724 11572 12733
rect 13820 12724 13872 12776
rect 14556 12767 14608 12776
rect 14556 12733 14565 12767
rect 14565 12733 14599 12767
rect 14599 12733 14608 12767
rect 14556 12724 14608 12733
rect 4068 12656 4120 12708
rect 16028 12631 16080 12640
rect 16028 12597 16037 12631
rect 16037 12597 16071 12631
rect 16071 12597 16080 12631
rect 16028 12588 16080 12597
rect 2985 12486 3037 12538
rect 3049 12486 3101 12538
rect 3113 12486 3165 12538
rect 3177 12486 3229 12538
rect 3241 12486 3293 12538
rect 7056 12486 7108 12538
rect 7120 12486 7172 12538
rect 7184 12486 7236 12538
rect 7248 12486 7300 12538
rect 7312 12486 7364 12538
rect 11127 12486 11179 12538
rect 11191 12486 11243 12538
rect 11255 12486 11307 12538
rect 11319 12486 11371 12538
rect 11383 12486 11435 12538
rect 15198 12486 15250 12538
rect 15262 12486 15314 12538
rect 15326 12486 15378 12538
rect 15390 12486 15442 12538
rect 15454 12486 15506 12538
rect 1676 12384 1728 12436
rect 3332 12384 3384 12436
rect 5540 12427 5592 12436
rect 5540 12393 5549 12427
rect 5549 12393 5583 12427
rect 5583 12393 5592 12427
rect 5540 12384 5592 12393
rect 7472 12427 7524 12436
rect 7472 12393 7481 12427
rect 7481 12393 7515 12427
rect 7515 12393 7524 12427
rect 7472 12384 7524 12393
rect 10876 12384 10928 12436
rect 12900 12384 12952 12436
rect 14556 12427 14608 12436
rect 14556 12393 14565 12427
rect 14565 12393 14599 12427
rect 14599 12393 14608 12427
rect 14556 12384 14608 12393
rect 16212 12427 16264 12436
rect 16212 12393 16221 12427
rect 16221 12393 16255 12427
rect 16255 12393 16264 12427
rect 16212 12384 16264 12393
rect 4068 12291 4120 12300
rect 4068 12257 4077 12291
rect 4077 12257 4111 12291
rect 4111 12257 4120 12291
rect 4068 12248 4120 12257
rect 7380 12248 7432 12300
rect 8116 12291 8168 12300
rect 8116 12257 8125 12291
rect 8125 12257 8159 12291
rect 8159 12257 8168 12291
rect 8116 12248 8168 12257
rect 2688 12180 2740 12232
rect 2872 12112 2924 12164
rect 3424 12180 3476 12232
rect 5172 12180 5224 12232
rect 8208 12180 8260 12232
rect 8944 12248 8996 12300
rect 8668 12180 8720 12232
rect 13544 12248 13596 12300
rect 13728 12180 13780 12232
rect 13820 12180 13872 12232
rect 15108 12180 15160 12232
rect 15752 12180 15804 12232
rect 16028 12180 16080 12232
rect 4344 12112 4396 12164
rect 15568 12112 15620 12164
rect 16212 12112 16264 12164
rect 8668 12087 8720 12096
rect 8668 12053 8677 12087
rect 8677 12053 8711 12087
rect 8711 12053 8720 12087
rect 8668 12044 8720 12053
rect 10232 12044 10284 12096
rect 11060 12044 11112 12096
rect 3645 11942 3697 11994
rect 3709 11942 3761 11994
rect 3773 11942 3825 11994
rect 3837 11942 3889 11994
rect 3901 11942 3953 11994
rect 7716 11942 7768 11994
rect 7780 11942 7832 11994
rect 7844 11942 7896 11994
rect 7908 11942 7960 11994
rect 7972 11942 8024 11994
rect 11787 11942 11839 11994
rect 11851 11942 11903 11994
rect 11915 11942 11967 11994
rect 11979 11942 12031 11994
rect 12043 11942 12095 11994
rect 15858 11942 15910 11994
rect 15922 11942 15974 11994
rect 15986 11942 16038 11994
rect 16050 11942 16102 11994
rect 16114 11942 16166 11994
rect 6000 11840 6052 11892
rect 6460 11840 6512 11892
rect 8668 11840 8720 11892
rect 10232 11883 10284 11892
rect 10232 11849 10241 11883
rect 10241 11849 10275 11883
rect 10275 11849 10284 11883
rect 10232 11840 10284 11849
rect 10324 11840 10376 11892
rect 9772 11772 9824 11824
rect 4712 11704 4764 11756
rect 5816 11704 5868 11756
rect 5908 11747 5960 11756
rect 5908 11713 5917 11747
rect 5917 11713 5951 11747
rect 5951 11713 5960 11747
rect 5908 11704 5960 11713
rect 6736 11704 6788 11756
rect 6920 11704 6972 11756
rect 8208 11704 8260 11756
rect 5356 11636 5408 11688
rect 7564 11679 7616 11688
rect 7564 11645 7573 11679
rect 7573 11645 7607 11679
rect 7607 11645 7616 11679
rect 7564 11636 7616 11645
rect 10324 11747 10376 11756
rect 10324 11713 10333 11747
rect 10333 11713 10367 11747
rect 10367 11713 10376 11747
rect 10324 11704 10376 11713
rect 10416 11747 10468 11756
rect 10416 11713 10425 11747
rect 10425 11713 10459 11747
rect 10459 11713 10468 11747
rect 10416 11704 10468 11713
rect 13084 11772 13136 11824
rect 13728 11772 13780 11824
rect 15108 11883 15160 11892
rect 15108 11849 15117 11883
rect 15117 11849 15151 11883
rect 15151 11849 15160 11883
rect 15108 11840 15160 11849
rect 15752 11772 15804 11824
rect 11520 11747 11572 11756
rect 11520 11713 11529 11747
rect 11529 11713 11563 11747
rect 11563 11713 11572 11747
rect 11520 11704 11572 11713
rect 10692 11636 10744 11688
rect 11796 11679 11848 11688
rect 11796 11645 11805 11679
rect 11805 11645 11839 11679
rect 11839 11645 11848 11679
rect 11796 11636 11848 11645
rect 13636 11679 13688 11688
rect 13636 11645 13645 11679
rect 13645 11645 13679 11679
rect 13679 11645 13688 11679
rect 13636 11636 13688 11645
rect 13728 11636 13780 11688
rect 14924 11704 14976 11756
rect 16488 11747 16540 11756
rect 16488 11713 16497 11747
rect 16497 11713 16531 11747
rect 16531 11713 16540 11747
rect 16488 11704 16540 11713
rect 16580 11704 16632 11756
rect 15568 11636 15620 11688
rect 16212 11679 16264 11688
rect 16212 11645 16221 11679
rect 16221 11645 16255 11679
rect 16255 11645 16264 11679
rect 16212 11636 16264 11645
rect 4252 11500 4304 11552
rect 6920 11500 6972 11552
rect 9772 11500 9824 11552
rect 10876 11500 10928 11552
rect 11520 11500 11572 11552
rect 13268 11543 13320 11552
rect 13268 11509 13277 11543
rect 13277 11509 13311 11543
rect 13311 11509 13320 11543
rect 13268 11500 13320 11509
rect 15108 11500 15160 11552
rect 15660 11500 15712 11552
rect 15752 11500 15804 11552
rect 2985 11398 3037 11450
rect 3049 11398 3101 11450
rect 3113 11398 3165 11450
rect 3177 11398 3229 11450
rect 3241 11398 3293 11450
rect 7056 11398 7108 11450
rect 7120 11398 7172 11450
rect 7184 11398 7236 11450
rect 7248 11398 7300 11450
rect 7312 11398 7364 11450
rect 11127 11398 11179 11450
rect 11191 11398 11243 11450
rect 11255 11398 11307 11450
rect 11319 11398 11371 11450
rect 11383 11398 11435 11450
rect 15198 11398 15250 11450
rect 15262 11398 15314 11450
rect 15326 11398 15378 11450
rect 15390 11398 15442 11450
rect 15454 11398 15506 11450
rect 2872 11296 2924 11348
rect 5816 11296 5868 11348
rect 10692 11339 10744 11348
rect 10692 11305 10701 11339
rect 10701 11305 10735 11339
rect 10735 11305 10744 11339
rect 10692 11296 10744 11305
rect 11796 11296 11848 11348
rect 13636 11296 13688 11348
rect 1400 11203 1452 11212
rect 1400 11169 1409 11203
rect 1409 11169 1443 11203
rect 1443 11169 1452 11203
rect 1400 11160 1452 11169
rect 6920 11228 6972 11280
rect 4252 11203 4304 11212
rect 4252 11169 4261 11203
rect 4261 11169 4295 11203
rect 4295 11169 4304 11203
rect 4252 11160 4304 11169
rect 4344 11160 4396 11212
rect 5172 11160 5224 11212
rect 2780 11092 2832 11144
rect 4160 11135 4212 11144
rect 4160 11101 4169 11135
rect 4169 11101 4203 11135
rect 4203 11101 4212 11135
rect 4160 11092 4212 11101
rect 4804 11067 4856 11076
rect 4804 11033 4813 11067
rect 4813 11033 4847 11067
rect 4847 11033 4856 11067
rect 4804 11024 4856 11033
rect 6828 11092 6880 11144
rect 8392 11160 8444 11212
rect 8668 11203 8720 11212
rect 8668 11169 8677 11203
rect 8677 11169 8711 11203
rect 8711 11169 8720 11203
rect 8668 11160 8720 11169
rect 9312 11160 9364 11212
rect 10876 11203 10928 11212
rect 10876 11169 10885 11203
rect 10885 11169 10919 11203
rect 10919 11169 10928 11203
rect 10876 11160 10928 11169
rect 12808 11203 12860 11212
rect 12808 11169 12817 11203
rect 12817 11169 12851 11203
rect 12851 11169 12860 11203
rect 12808 11160 12860 11169
rect 14280 11160 14332 11212
rect 15660 11160 15712 11212
rect 16488 11160 16540 11212
rect 10968 11135 11020 11144
rect 10968 11101 10977 11135
rect 10977 11101 11011 11135
rect 11011 11101 11020 11135
rect 10968 11092 11020 11101
rect 12440 11092 12492 11144
rect 13268 11092 13320 11144
rect 17040 11135 17092 11144
rect 17040 11101 17049 11135
rect 17049 11101 17083 11135
rect 17083 11101 17092 11135
rect 17040 11092 17092 11101
rect 1400 10956 1452 11008
rect 2596 10956 2648 11008
rect 9220 11067 9272 11076
rect 9220 11033 9229 11067
rect 9229 11033 9263 11067
rect 9263 11033 9272 11067
rect 9220 11024 9272 11033
rect 10784 11024 10836 11076
rect 15752 11024 15804 11076
rect 8484 10956 8536 11008
rect 16580 10956 16632 11008
rect 16856 10999 16908 11008
rect 16856 10965 16865 10999
rect 16865 10965 16899 10999
rect 16899 10965 16908 10999
rect 16856 10956 16908 10965
rect 3645 10854 3697 10906
rect 3709 10854 3761 10906
rect 3773 10854 3825 10906
rect 3837 10854 3889 10906
rect 3901 10854 3953 10906
rect 7716 10854 7768 10906
rect 7780 10854 7832 10906
rect 7844 10854 7896 10906
rect 7908 10854 7960 10906
rect 7972 10854 8024 10906
rect 11787 10854 11839 10906
rect 11851 10854 11903 10906
rect 11915 10854 11967 10906
rect 11979 10854 12031 10906
rect 12043 10854 12095 10906
rect 15858 10854 15910 10906
rect 15922 10854 15974 10906
rect 15986 10854 16038 10906
rect 16050 10854 16102 10906
rect 16114 10854 16166 10906
rect 2780 10752 2832 10804
rect 848 10616 900 10668
rect 2044 10616 2096 10668
rect 4160 10752 4212 10804
rect 2596 10659 2648 10668
rect 2596 10625 2605 10659
rect 2605 10625 2639 10659
rect 2639 10625 2648 10659
rect 2596 10616 2648 10625
rect 4804 10752 4856 10804
rect 5356 10752 5408 10804
rect 6736 10752 6788 10804
rect 5816 10659 5868 10668
rect 5816 10625 5825 10659
rect 5825 10625 5859 10659
rect 5859 10625 5868 10659
rect 5816 10616 5868 10625
rect 4712 10548 4764 10600
rect 5908 10480 5960 10532
rect 7564 10616 7616 10668
rect 8392 10752 8444 10804
rect 9220 10752 9272 10804
rect 10416 10795 10468 10804
rect 10416 10761 10425 10795
rect 10425 10761 10459 10795
rect 10459 10761 10468 10795
rect 10416 10752 10468 10761
rect 12808 10752 12860 10804
rect 14924 10752 14976 10804
rect 16212 10795 16264 10804
rect 16212 10761 16221 10795
rect 16221 10761 16255 10795
rect 16255 10761 16264 10795
rect 16212 10752 16264 10761
rect 8484 10684 8536 10736
rect 8760 10616 8812 10668
rect 9772 10659 9824 10668
rect 9772 10625 9781 10659
rect 9781 10625 9815 10659
rect 9815 10625 9824 10659
rect 9772 10616 9824 10625
rect 10692 10684 10744 10736
rect 10416 10659 10468 10668
rect 10416 10625 10425 10659
rect 10425 10625 10459 10659
rect 10459 10625 10468 10659
rect 10416 10616 10468 10625
rect 12440 10659 12492 10668
rect 12440 10625 12449 10659
rect 12449 10625 12483 10659
rect 12483 10625 12492 10659
rect 12440 10616 12492 10625
rect 15200 10684 15252 10736
rect 13268 10616 13320 10668
rect 16580 10752 16632 10804
rect 16488 10727 16540 10736
rect 16488 10693 16497 10727
rect 16497 10693 16531 10727
rect 16531 10693 16540 10727
rect 16488 10684 16540 10693
rect 12808 10591 12860 10600
rect 12808 10557 12817 10591
rect 12817 10557 12851 10591
rect 12851 10557 12860 10591
rect 12808 10548 12860 10557
rect 14924 10548 14976 10600
rect 16856 10616 16908 10668
rect 17040 10659 17092 10668
rect 17040 10625 17049 10659
rect 17049 10625 17083 10659
rect 17083 10625 17092 10659
rect 17040 10616 17092 10625
rect 16948 10548 17000 10600
rect 10968 10480 11020 10532
rect 2872 10412 2924 10464
rect 8208 10412 8260 10464
rect 11704 10412 11756 10464
rect 13728 10412 13780 10464
rect 2985 10310 3037 10362
rect 3049 10310 3101 10362
rect 3113 10310 3165 10362
rect 3177 10310 3229 10362
rect 3241 10310 3293 10362
rect 7056 10310 7108 10362
rect 7120 10310 7172 10362
rect 7184 10310 7236 10362
rect 7248 10310 7300 10362
rect 7312 10310 7364 10362
rect 11127 10310 11179 10362
rect 11191 10310 11243 10362
rect 11255 10310 11307 10362
rect 11319 10310 11371 10362
rect 11383 10310 11435 10362
rect 15198 10310 15250 10362
rect 15262 10310 15314 10362
rect 15326 10310 15378 10362
rect 15390 10310 15442 10362
rect 15454 10310 15506 10362
rect 13268 10251 13320 10260
rect 13268 10217 13277 10251
rect 13277 10217 13311 10251
rect 13311 10217 13320 10251
rect 13268 10208 13320 10217
rect 14924 10208 14976 10260
rect 15568 10208 15620 10260
rect 11704 10115 11756 10124
rect 11704 10081 11713 10115
rect 11713 10081 11747 10115
rect 11747 10081 11756 10115
rect 11704 10072 11756 10081
rect 13084 10072 13136 10124
rect 1400 10047 1452 10056
rect 1400 10013 1409 10047
rect 1409 10013 1443 10047
rect 1443 10013 1452 10047
rect 1400 10004 1452 10013
rect 8116 10004 8168 10056
rect 8300 10004 8352 10056
rect 11428 10047 11480 10056
rect 11428 10013 11437 10047
rect 11437 10013 11471 10047
rect 11471 10013 11480 10047
rect 11428 10004 11480 10013
rect 15384 10115 15436 10124
rect 15384 10081 15393 10115
rect 15393 10081 15427 10115
rect 15427 10081 15436 10115
rect 15384 10072 15436 10081
rect 13728 10047 13780 10056
rect 13728 10013 13737 10047
rect 13737 10013 13771 10047
rect 13771 10013 13780 10047
rect 13728 10004 13780 10013
rect 15752 10004 15804 10056
rect 16488 10004 16540 10056
rect 16856 10004 16908 10056
rect 12440 9936 12492 9988
rect 2964 9868 3016 9920
rect 8484 9868 8536 9920
rect 12716 9868 12768 9920
rect 16212 9868 16264 9920
rect 3645 9766 3697 9818
rect 3709 9766 3761 9818
rect 3773 9766 3825 9818
rect 3837 9766 3889 9818
rect 3901 9766 3953 9818
rect 7716 9766 7768 9818
rect 7780 9766 7832 9818
rect 7844 9766 7896 9818
rect 7908 9766 7960 9818
rect 7972 9766 8024 9818
rect 11787 9766 11839 9818
rect 11851 9766 11903 9818
rect 11915 9766 11967 9818
rect 11979 9766 12031 9818
rect 12043 9766 12095 9818
rect 15858 9766 15910 9818
rect 15922 9766 15974 9818
rect 15986 9766 16038 9818
rect 16050 9766 16102 9818
rect 16114 9766 16166 9818
rect 2872 9664 2924 9716
rect 12808 9707 12860 9716
rect 12808 9673 12817 9707
rect 12817 9673 12851 9707
rect 12851 9673 12860 9707
rect 12808 9664 12860 9673
rect 15384 9664 15436 9716
rect 16212 9664 16264 9716
rect 1584 9639 1636 9648
rect 1584 9605 1593 9639
rect 1593 9605 1627 9639
rect 1627 9605 1636 9639
rect 1584 9596 1636 9605
rect 3516 9596 3568 9648
rect 3976 9596 4028 9648
rect 8208 9596 8260 9648
rect 9956 9596 10008 9648
rect 13084 9639 13136 9648
rect 13084 9605 13093 9639
rect 13093 9605 13127 9639
rect 13127 9605 13136 9639
rect 13084 9596 13136 9605
rect 2044 9503 2096 9512
rect 2044 9469 2053 9503
rect 2053 9469 2087 9503
rect 2087 9469 2096 9503
rect 2044 9460 2096 9469
rect 2412 9503 2464 9512
rect 2412 9469 2421 9503
rect 2421 9469 2455 9503
rect 2455 9469 2464 9503
rect 2412 9460 2464 9469
rect 2688 9571 2740 9580
rect 2688 9537 2697 9571
rect 2697 9537 2731 9571
rect 2731 9537 2740 9571
rect 2688 9528 2740 9537
rect 2872 9571 2924 9580
rect 2872 9537 2881 9571
rect 2881 9537 2915 9571
rect 2915 9537 2924 9571
rect 2872 9528 2924 9537
rect 2964 9571 3016 9580
rect 2964 9537 2973 9571
rect 2973 9537 3007 9571
rect 3007 9537 3016 9571
rect 2964 9528 3016 9537
rect 1584 9392 1636 9444
rect 3332 9528 3384 9580
rect 5724 9571 5776 9580
rect 5724 9537 5733 9571
rect 5733 9537 5767 9571
rect 5767 9537 5776 9571
rect 5724 9528 5776 9537
rect 5816 9571 5868 9580
rect 5816 9537 5825 9571
rect 5825 9537 5859 9571
rect 5859 9537 5868 9571
rect 5816 9528 5868 9537
rect 5540 9460 5592 9512
rect 8116 9528 8168 9580
rect 7380 9460 7432 9512
rect 8668 9528 8720 9580
rect 12808 9571 12860 9580
rect 12808 9537 12817 9571
rect 12817 9537 12851 9571
rect 12851 9537 12860 9571
rect 12808 9528 12860 9537
rect 13728 9528 13780 9580
rect 8300 9503 8352 9512
rect 8300 9469 8309 9503
rect 8309 9469 8343 9503
rect 8343 9469 8352 9503
rect 8300 9460 8352 9469
rect 8484 9503 8536 9512
rect 8484 9469 8493 9503
rect 8493 9469 8527 9503
rect 8527 9469 8536 9503
rect 8484 9460 8536 9469
rect 9128 9503 9180 9512
rect 9128 9469 9137 9503
rect 9137 9469 9171 9503
rect 9171 9469 9180 9503
rect 9128 9460 9180 9469
rect 1492 9367 1544 9376
rect 1492 9333 1501 9367
rect 1501 9333 1535 9367
rect 1535 9333 1544 9367
rect 1492 9324 1544 9333
rect 1676 9324 1728 9376
rect 8852 9392 8904 9444
rect 15936 9528 15988 9580
rect 16304 9528 16356 9580
rect 16856 9528 16908 9580
rect 16120 9460 16172 9512
rect 6368 9324 6420 9376
rect 6920 9324 6972 9376
rect 10692 9324 10744 9376
rect 2985 9222 3037 9274
rect 3049 9222 3101 9274
rect 3113 9222 3165 9274
rect 3177 9222 3229 9274
rect 3241 9222 3293 9274
rect 7056 9222 7108 9274
rect 7120 9222 7172 9274
rect 7184 9222 7236 9274
rect 7248 9222 7300 9274
rect 7312 9222 7364 9274
rect 11127 9222 11179 9274
rect 11191 9222 11243 9274
rect 11255 9222 11307 9274
rect 11319 9222 11371 9274
rect 11383 9222 11435 9274
rect 15198 9222 15250 9274
rect 15262 9222 15314 9274
rect 15326 9222 15378 9274
rect 15390 9222 15442 9274
rect 15454 9222 15506 9274
rect 2688 9120 2740 9172
rect 1676 9027 1728 9036
rect 1676 8993 1685 9027
rect 1685 8993 1719 9027
rect 1719 8993 1728 9027
rect 1676 8984 1728 8993
rect 3332 9163 3384 9172
rect 3332 9129 3341 9163
rect 3341 9129 3375 9163
rect 3375 9129 3384 9163
rect 3332 9120 3384 9129
rect 7380 9120 7432 9172
rect 8300 9120 8352 9172
rect 15752 9120 15804 9172
rect 9128 9052 9180 9104
rect 15936 9120 15988 9172
rect 6920 9027 6972 9036
rect 6920 8993 6929 9027
rect 6929 8993 6963 9027
rect 6963 8993 6972 9027
rect 6920 8984 6972 8993
rect 10600 9027 10652 9036
rect 10600 8993 10609 9027
rect 10609 8993 10643 9027
rect 10643 8993 10652 9027
rect 10600 8984 10652 8993
rect 16120 9027 16172 9036
rect 16120 8993 16129 9027
rect 16129 8993 16163 9027
rect 16163 8993 16172 9027
rect 16120 8984 16172 8993
rect 3424 8959 3476 8968
rect 3424 8925 3433 8959
rect 3433 8925 3467 8959
rect 3467 8925 3476 8959
rect 3424 8916 3476 8925
rect 3516 8959 3568 8968
rect 3516 8925 3525 8959
rect 3525 8925 3559 8959
rect 3559 8925 3568 8959
rect 3516 8916 3568 8925
rect 3700 8848 3752 8900
rect 1584 8780 1636 8832
rect 6184 8916 6236 8968
rect 6368 8959 6420 8968
rect 6368 8925 6377 8959
rect 6377 8925 6411 8959
rect 6411 8925 6420 8959
rect 6368 8916 6420 8925
rect 6552 8959 6604 8968
rect 6552 8925 6561 8959
rect 6561 8925 6595 8959
rect 6595 8925 6604 8959
rect 6552 8916 6604 8925
rect 8760 8959 8812 8968
rect 8760 8925 8769 8959
rect 8769 8925 8803 8959
rect 8803 8925 8812 8959
rect 8760 8916 8812 8925
rect 8852 8916 8904 8968
rect 5356 8848 5408 8900
rect 7380 8848 7432 8900
rect 4712 8780 4764 8832
rect 5540 8823 5592 8832
rect 5540 8789 5549 8823
rect 5549 8789 5583 8823
rect 5583 8789 5592 8823
rect 5540 8780 5592 8789
rect 6460 8823 6512 8832
rect 6460 8789 6469 8823
rect 6469 8789 6503 8823
rect 6503 8789 6512 8823
rect 6460 8780 6512 8789
rect 8392 8823 8444 8832
rect 8392 8789 8401 8823
rect 8401 8789 8435 8823
rect 8435 8789 8444 8823
rect 8668 8891 8720 8900
rect 8668 8857 8677 8891
rect 8677 8857 8711 8891
rect 8711 8857 8720 8891
rect 8668 8848 8720 8857
rect 10692 8959 10744 8968
rect 10692 8925 10701 8959
rect 10701 8925 10735 8959
rect 10735 8925 10744 8959
rect 10692 8916 10744 8925
rect 14096 8959 14148 8968
rect 14096 8925 14105 8959
rect 14105 8925 14139 8959
rect 14139 8925 14148 8959
rect 14096 8916 14148 8925
rect 13912 8848 13964 8900
rect 8392 8780 8444 8789
rect 11060 8823 11112 8832
rect 11060 8789 11069 8823
rect 11069 8789 11103 8823
rect 11103 8789 11112 8823
rect 11060 8780 11112 8789
rect 15016 8780 15068 8832
rect 16304 8916 16356 8968
rect 16856 8959 16908 8968
rect 16856 8925 16865 8959
rect 16865 8925 16899 8959
rect 16899 8925 16908 8959
rect 16856 8916 16908 8925
rect 16948 8959 17000 8968
rect 16948 8925 16957 8959
rect 16957 8925 16991 8959
rect 16991 8925 17000 8959
rect 16948 8916 17000 8925
rect 16396 8848 16448 8900
rect 3645 8678 3697 8730
rect 3709 8678 3761 8730
rect 3773 8678 3825 8730
rect 3837 8678 3889 8730
rect 3901 8678 3953 8730
rect 7716 8678 7768 8730
rect 7780 8678 7832 8730
rect 7844 8678 7896 8730
rect 7908 8678 7960 8730
rect 7972 8678 8024 8730
rect 11787 8678 11839 8730
rect 11851 8678 11903 8730
rect 11915 8678 11967 8730
rect 11979 8678 12031 8730
rect 12043 8678 12095 8730
rect 15858 8678 15910 8730
rect 15922 8678 15974 8730
rect 15986 8678 16038 8730
rect 16050 8678 16102 8730
rect 16114 8678 16166 8730
rect 2044 8576 2096 8628
rect 5724 8576 5776 8628
rect 3976 8508 4028 8560
rect 848 8440 900 8492
rect 1676 8483 1728 8492
rect 1676 8449 1685 8483
rect 1685 8449 1719 8483
rect 1719 8449 1728 8483
rect 1676 8440 1728 8449
rect 4712 8483 4764 8492
rect 4712 8449 4721 8483
rect 4721 8449 4755 8483
rect 4755 8449 4764 8483
rect 4712 8440 4764 8449
rect 2412 8236 2464 8288
rect 3424 8236 3476 8288
rect 3976 8236 4028 8288
rect 5264 8236 5316 8288
rect 5540 8508 5592 8560
rect 6184 8440 6236 8492
rect 6552 8619 6604 8628
rect 6552 8585 6561 8619
rect 6561 8585 6595 8619
rect 6595 8585 6604 8619
rect 6552 8576 6604 8585
rect 8116 8576 8168 8628
rect 10600 8619 10652 8628
rect 10600 8585 10609 8619
rect 10609 8585 10643 8619
rect 10643 8585 10652 8619
rect 10600 8576 10652 8585
rect 10692 8576 10744 8628
rect 13912 8619 13964 8628
rect 13912 8585 13921 8619
rect 13921 8585 13955 8619
rect 13955 8585 13964 8619
rect 13912 8576 13964 8585
rect 16304 8576 16356 8628
rect 16856 8619 16908 8628
rect 16856 8585 16865 8619
rect 16865 8585 16899 8619
rect 16899 8585 16908 8619
rect 16856 8576 16908 8585
rect 6736 8440 6788 8492
rect 8392 8508 8444 8560
rect 6460 8372 6512 8424
rect 6920 8372 6972 8424
rect 7564 8372 7616 8424
rect 8668 8440 8720 8492
rect 11060 8508 11112 8560
rect 12440 8508 12492 8560
rect 15016 8551 15068 8560
rect 15016 8517 15025 8551
rect 15025 8517 15059 8551
rect 15059 8517 15068 8551
rect 15016 8508 15068 8517
rect 16396 8508 16448 8560
rect 10416 8415 10468 8424
rect 10416 8381 10425 8415
rect 10425 8381 10459 8415
rect 10459 8381 10468 8415
rect 10416 8372 10468 8381
rect 11520 8415 11572 8424
rect 11520 8381 11529 8415
rect 11529 8381 11563 8415
rect 11563 8381 11572 8415
rect 11520 8372 11572 8381
rect 13636 8440 13688 8492
rect 14096 8440 14148 8492
rect 14556 8440 14608 8492
rect 17040 8483 17092 8492
rect 17040 8449 17049 8483
rect 17049 8449 17083 8483
rect 17083 8449 17092 8483
rect 17040 8440 17092 8449
rect 13452 8415 13504 8424
rect 13452 8381 13461 8415
rect 13461 8381 13495 8415
rect 13495 8381 13504 8415
rect 13452 8372 13504 8381
rect 10784 8304 10836 8356
rect 9772 8279 9824 8288
rect 9772 8245 9781 8279
rect 9781 8245 9815 8279
rect 9815 8245 9824 8279
rect 9772 8236 9824 8245
rect 2985 8134 3037 8186
rect 3049 8134 3101 8186
rect 3113 8134 3165 8186
rect 3177 8134 3229 8186
rect 3241 8134 3293 8186
rect 7056 8134 7108 8186
rect 7120 8134 7172 8186
rect 7184 8134 7236 8186
rect 7248 8134 7300 8186
rect 7312 8134 7364 8186
rect 11127 8134 11179 8186
rect 11191 8134 11243 8186
rect 11255 8134 11307 8186
rect 11319 8134 11371 8186
rect 11383 8134 11435 8186
rect 15198 8134 15250 8186
rect 15262 8134 15314 8186
rect 15326 8134 15378 8186
rect 15390 8134 15442 8186
rect 15454 8134 15506 8186
rect 2228 8032 2280 8084
rect 10784 8075 10836 8084
rect 10784 8041 10793 8075
rect 10793 8041 10827 8075
rect 10827 8041 10836 8075
rect 10784 8032 10836 8041
rect 13452 8032 13504 8084
rect 848 7828 900 7880
rect 8208 7964 8260 8016
rect 8668 7964 8720 8016
rect 8300 7896 8352 7948
rect 9772 7896 9824 7948
rect 6920 7760 6972 7812
rect 3148 7735 3200 7744
rect 3148 7701 3157 7735
rect 3157 7701 3191 7735
rect 3191 7701 3200 7735
rect 3148 7692 3200 7701
rect 3424 7692 3476 7744
rect 7564 7692 7616 7744
rect 8208 7871 8260 7880
rect 8208 7837 8217 7871
rect 8217 7837 8251 7871
rect 8251 7837 8260 7871
rect 8208 7828 8260 7837
rect 8116 7760 8168 7812
rect 9128 7760 9180 7812
rect 9956 7760 10008 7812
rect 10876 7760 10928 7812
rect 13544 7828 13596 7880
rect 17040 7871 17092 7880
rect 17040 7837 17049 7871
rect 17049 7837 17083 7871
rect 17083 7837 17092 7871
rect 17040 7828 17092 7837
rect 14004 7760 14056 7812
rect 8484 7692 8536 7744
rect 10692 7735 10744 7744
rect 10692 7701 10701 7735
rect 10701 7701 10735 7735
rect 10735 7701 10744 7735
rect 10692 7692 10744 7701
rect 12716 7692 12768 7744
rect 14280 7692 14332 7744
rect 3645 7590 3697 7642
rect 3709 7590 3761 7642
rect 3773 7590 3825 7642
rect 3837 7590 3889 7642
rect 3901 7590 3953 7642
rect 7716 7590 7768 7642
rect 7780 7590 7832 7642
rect 7844 7590 7896 7642
rect 7908 7590 7960 7642
rect 7972 7590 8024 7642
rect 11787 7590 11839 7642
rect 11851 7590 11903 7642
rect 11915 7590 11967 7642
rect 11979 7590 12031 7642
rect 12043 7590 12095 7642
rect 15858 7590 15910 7642
rect 15922 7590 15974 7642
rect 15986 7590 16038 7642
rect 16050 7590 16102 7642
rect 16114 7590 16166 7642
rect 6184 7531 6236 7540
rect 6184 7497 6193 7531
rect 6193 7497 6227 7531
rect 6227 7497 6236 7531
rect 6184 7488 6236 7497
rect 7380 7488 7432 7540
rect 7656 7488 7708 7540
rect 8116 7531 8168 7540
rect 8116 7497 8125 7531
rect 8125 7497 8159 7531
rect 8159 7497 8168 7531
rect 8116 7488 8168 7497
rect 10416 7488 10468 7540
rect 3608 7420 3660 7472
rect 3976 7420 4028 7472
rect 2228 7395 2280 7404
rect 2228 7361 2237 7395
rect 2237 7361 2271 7395
rect 2271 7361 2280 7395
rect 2228 7352 2280 7361
rect 2412 7352 2464 7404
rect 4712 7420 4764 7472
rect 5264 7420 5316 7472
rect 6920 7420 6972 7472
rect 7288 7420 7340 7472
rect 10692 7420 10744 7472
rect 12440 7420 12492 7472
rect 14004 7531 14056 7540
rect 14004 7497 14013 7531
rect 14013 7497 14047 7531
rect 14047 7497 14056 7531
rect 14004 7488 14056 7497
rect 13452 7420 13504 7472
rect 14280 7463 14332 7472
rect 14280 7429 14289 7463
rect 14289 7429 14323 7463
rect 14323 7429 14332 7463
rect 14280 7420 14332 7429
rect 16396 7420 16448 7472
rect 8024 7352 8076 7404
rect 8668 7352 8720 7404
rect 10324 7352 10376 7404
rect 10876 7352 10928 7404
rect 13636 7395 13688 7404
rect 13636 7361 13645 7395
rect 13645 7361 13679 7395
rect 13679 7361 13688 7395
rect 13636 7352 13688 7361
rect 13820 7352 13872 7404
rect 14556 7395 14608 7404
rect 14556 7361 14565 7395
rect 14565 7361 14599 7395
rect 14599 7361 14608 7395
rect 14556 7352 14608 7361
rect 17040 7395 17092 7404
rect 17040 7361 17049 7395
rect 17049 7361 17083 7395
rect 17083 7361 17092 7395
rect 17040 7352 17092 7361
rect 3424 7284 3476 7336
rect 4068 7327 4120 7336
rect 4068 7293 4077 7327
rect 4077 7293 4111 7327
rect 4111 7293 4120 7327
rect 4068 7284 4120 7293
rect 2872 7148 2924 7200
rect 3976 7148 4028 7200
rect 7380 7284 7432 7336
rect 8484 7327 8536 7336
rect 8484 7293 8493 7327
rect 8493 7293 8527 7327
rect 8527 7293 8536 7327
rect 8484 7284 8536 7293
rect 9128 7284 9180 7336
rect 11520 7327 11572 7336
rect 11520 7293 11529 7327
rect 11529 7293 11563 7327
rect 11563 7293 11572 7327
rect 11520 7284 11572 7293
rect 13544 7327 13596 7336
rect 13544 7293 13553 7327
rect 13553 7293 13587 7327
rect 13587 7293 13596 7327
rect 13544 7284 13596 7293
rect 15568 7284 15620 7336
rect 16304 7191 16356 7200
rect 16304 7157 16313 7191
rect 16313 7157 16347 7191
rect 16347 7157 16356 7191
rect 16304 7148 16356 7157
rect 16672 7148 16724 7200
rect 2985 7046 3037 7098
rect 3049 7046 3101 7098
rect 3113 7046 3165 7098
rect 3177 7046 3229 7098
rect 3241 7046 3293 7098
rect 7056 7046 7108 7098
rect 7120 7046 7172 7098
rect 7184 7046 7236 7098
rect 7248 7046 7300 7098
rect 7312 7046 7364 7098
rect 11127 7046 11179 7098
rect 11191 7046 11243 7098
rect 11255 7046 11307 7098
rect 11319 7046 11371 7098
rect 11383 7046 11435 7098
rect 15198 7046 15250 7098
rect 15262 7046 15314 7098
rect 15326 7046 15378 7098
rect 15390 7046 15442 7098
rect 15454 7046 15506 7098
rect 3332 6740 3384 6792
rect 4068 6944 4120 6996
rect 8208 6944 8260 6996
rect 13544 6944 13596 6996
rect 6920 6808 6972 6860
rect 7564 6808 7616 6860
rect 15568 6808 15620 6860
rect 16212 6808 16264 6860
rect 3976 6783 4028 6792
rect 3976 6749 3985 6783
rect 3985 6749 4019 6783
rect 4019 6749 4028 6783
rect 3976 6740 4028 6749
rect 4068 6740 4120 6792
rect 1584 6672 1636 6724
rect 3608 6672 3660 6724
rect 3424 6604 3476 6656
rect 5080 6647 5132 6656
rect 5080 6613 5089 6647
rect 5089 6613 5123 6647
rect 5123 6613 5132 6647
rect 5080 6604 5132 6613
rect 6920 6672 6972 6724
rect 5816 6604 5868 6656
rect 6460 6647 6512 6656
rect 6460 6613 6469 6647
rect 6469 6613 6503 6647
rect 6503 6613 6512 6647
rect 6460 6604 6512 6613
rect 8116 6740 8168 6792
rect 8300 6783 8352 6792
rect 8300 6749 8309 6783
rect 8309 6749 8343 6783
rect 8343 6749 8352 6783
rect 8300 6740 8352 6749
rect 13452 6740 13504 6792
rect 13728 6740 13780 6792
rect 14280 6740 14332 6792
rect 10968 6672 11020 6724
rect 12808 6672 12860 6724
rect 15660 6740 15712 6792
rect 16304 6740 16356 6792
rect 16672 6783 16724 6792
rect 16672 6749 16681 6783
rect 16681 6749 16715 6783
rect 16715 6749 16724 6783
rect 16672 6740 16724 6749
rect 16856 6740 16908 6792
rect 15752 6672 15804 6724
rect 8116 6604 8168 6656
rect 10048 6604 10100 6656
rect 12716 6604 12768 6656
rect 16120 6604 16172 6656
rect 16304 6647 16356 6656
rect 16304 6613 16313 6647
rect 16313 6613 16347 6647
rect 16347 6613 16356 6647
rect 16304 6604 16356 6613
rect 3645 6502 3697 6554
rect 3709 6502 3761 6554
rect 3773 6502 3825 6554
rect 3837 6502 3889 6554
rect 3901 6502 3953 6554
rect 7716 6502 7768 6554
rect 7780 6502 7832 6554
rect 7844 6502 7896 6554
rect 7908 6502 7960 6554
rect 7972 6502 8024 6554
rect 11787 6502 11839 6554
rect 11851 6502 11903 6554
rect 11915 6502 11967 6554
rect 11979 6502 12031 6554
rect 12043 6502 12095 6554
rect 15858 6502 15910 6554
rect 15922 6502 15974 6554
rect 15986 6502 16038 6554
rect 16050 6502 16102 6554
rect 16114 6502 16166 6554
rect 2780 6400 2832 6452
rect 5080 6400 5132 6452
rect 6460 6400 6512 6452
rect 14464 6400 14516 6452
rect 9956 6332 10008 6384
rect 10968 6332 11020 6384
rect 2504 6264 2556 6316
rect 2872 6196 2924 6248
rect 8208 6264 8260 6316
rect 9128 6264 9180 6316
rect 9864 6196 9916 6248
rect 13728 6307 13780 6316
rect 13728 6273 13737 6307
rect 13737 6273 13771 6307
rect 13771 6273 13780 6307
rect 13728 6264 13780 6273
rect 13912 6264 13964 6316
rect 15752 6307 15804 6316
rect 15752 6273 15761 6307
rect 15761 6273 15795 6307
rect 15795 6273 15804 6307
rect 15752 6264 15804 6273
rect 16212 6264 16264 6316
rect 14556 6196 14608 6248
rect 10784 6128 10836 6180
rect 11704 6128 11756 6180
rect 3332 6060 3384 6112
rect 10048 6060 10100 6112
rect 10600 6060 10652 6112
rect 14004 6060 14056 6112
rect 15752 6060 15804 6112
rect 2985 5958 3037 6010
rect 3049 5958 3101 6010
rect 3113 5958 3165 6010
rect 3177 5958 3229 6010
rect 3241 5958 3293 6010
rect 7056 5958 7108 6010
rect 7120 5958 7172 6010
rect 7184 5958 7236 6010
rect 7248 5958 7300 6010
rect 7312 5958 7364 6010
rect 11127 5958 11179 6010
rect 11191 5958 11243 6010
rect 11255 5958 11307 6010
rect 11319 5958 11371 6010
rect 11383 5958 11435 6010
rect 15198 5958 15250 6010
rect 15262 5958 15314 6010
rect 15326 5958 15378 6010
rect 15390 5958 15442 6010
rect 15454 5958 15506 6010
rect 3148 5856 3200 5908
rect 3516 5856 3568 5908
rect 6920 5856 6972 5908
rect 7196 5856 7248 5908
rect 8208 5856 8260 5908
rect 9864 5899 9916 5908
rect 9864 5865 9873 5899
rect 9873 5865 9907 5899
rect 9907 5865 9916 5899
rect 9864 5856 9916 5865
rect 9956 5856 10008 5908
rect 12440 5856 12492 5908
rect 13912 5899 13964 5908
rect 13912 5865 13921 5899
rect 13921 5865 13955 5899
rect 13955 5865 13964 5899
rect 13912 5856 13964 5865
rect 2504 5788 2556 5840
rect 7012 5788 7064 5840
rect 10692 5788 10744 5840
rect 10968 5788 11020 5840
rect 3332 5720 3384 5772
rect 3424 5763 3476 5772
rect 3424 5729 3433 5763
rect 3433 5729 3467 5763
rect 3467 5729 3476 5763
rect 3424 5720 3476 5729
rect 3516 5720 3568 5772
rect 6828 5720 6880 5772
rect 1400 5695 1452 5704
rect 1400 5661 1409 5695
rect 1409 5661 1443 5695
rect 1443 5661 1452 5695
rect 1400 5652 1452 5661
rect 2412 5695 2464 5704
rect 2412 5661 2421 5695
rect 2421 5661 2455 5695
rect 2455 5661 2464 5695
rect 2412 5652 2464 5661
rect 2504 5695 2556 5704
rect 2504 5661 2513 5695
rect 2513 5661 2547 5695
rect 2547 5661 2556 5695
rect 2504 5652 2556 5661
rect 2780 5652 2832 5704
rect 6920 5695 6972 5704
rect 6920 5661 6929 5695
rect 6929 5661 6963 5695
rect 6963 5661 6972 5695
rect 6920 5652 6972 5661
rect 7196 5695 7248 5704
rect 7196 5661 7205 5695
rect 7205 5661 7239 5695
rect 7239 5661 7248 5695
rect 7196 5652 7248 5661
rect 8208 5652 8260 5704
rect 10140 5695 10192 5704
rect 10140 5661 10149 5695
rect 10149 5661 10183 5695
rect 10183 5661 10192 5695
rect 10140 5652 10192 5661
rect 11520 5720 11572 5772
rect 10600 5695 10652 5704
rect 10600 5661 10609 5695
rect 10609 5661 10643 5695
rect 10643 5661 10652 5695
rect 10600 5652 10652 5661
rect 10784 5695 10836 5704
rect 10784 5661 10793 5695
rect 10793 5661 10827 5695
rect 10827 5661 10836 5695
rect 10784 5652 10836 5661
rect 14556 5788 14608 5840
rect 14464 5695 14516 5704
rect 14464 5661 14473 5695
rect 14473 5661 14507 5695
rect 14507 5661 14516 5695
rect 14464 5652 14516 5661
rect 15752 5763 15804 5772
rect 15752 5729 15761 5763
rect 15761 5729 15795 5763
rect 15795 5729 15804 5763
rect 15752 5720 15804 5729
rect 15660 5695 15712 5704
rect 15660 5661 15669 5695
rect 15669 5661 15703 5695
rect 15703 5661 15712 5695
rect 15660 5652 15712 5661
rect 17040 5695 17092 5704
rect 17040 5661 17049 5695
rect 17049 5661 17083 5695
rect 17083 5661 17092 5695
rect 17040 5652 17092 5661
rect 2872 5584 2924 5636
rect 3240 5584 3292 5636
rect 5080 5584 5132 5636
rect 2780 5559 2832 5568
rect 2780 5525 2789 5559
rect 2789 5525 2823 5559
rect 2823 5525 2832 5559
rect 2780 5516 2832 5525
rect 4528 5516 4580 5568
rect 6552 5516 6604 5568
rect 12440 5627 12492 5636
rect 12440 5593 12449 5627
rect 12449 5593 12483 5627
rect 12483 5593 12492 5627
rect 12440 5584 12492 5593
rect 12532 5584 12584 5636
rect 12900 5584 12952 5636
rect 10600 5559 10652 5568
rect 10600 5525 10609 5559
rect 10609 5525 10643 5559
rect 10643 5525 10652 5559
rect 10600 5516 10652 5525
rect 14096 5559 14148 5568
rect 14096 5525 14105 5559
rect 14105 5525 14139 5559
rect 14139 5525 14148 5559
rect 14096 5516 14148 5525
rect 16764 5516 16816 5568
rect 3645 5414 3697 5466
rect 3709 5414 3761 5466
rect 3773 5414 3825 5466
rect 3837 5414 3889 5466
rect 3901 5414 3953 5466
rect 7716 5414 7768 5466
rect 7780 5414 7832 5466
rect 7844 5414 7896 5466
rect 7908 5414 7960 5466
rect 7972 5414 8024 5466
rect 11787 5414 11839 5466
rect 11851 5414 11903 5466
rect 11915 5414 11967 5466
rect 11979 5414 12031 5466
rect 12043 5414 12095 5466
rect 15858 5414 15910 5466
rect 15922 5414 15974 5466
rect 15986 5414 16038 5466
rect 16050 5414 16102 5466
rect 16114 5414 16166 5466
rect 2780 5312 2832 5364
rect 3516 5355 3568 5364
rect 3516 5321 3525 5355
rect 3525 5321 3559 5355
rect 3559 5321 3568 5355
rect 3516 5312 3568 5321
rect 7012 5355 7064 5364
rect 7012 5321 7021 5355
rect 7021 5321 7055 5355
rect 7055 5321 7064 5355
rect 7012 5312 7064 5321
rect 7380 5312 7432 5364
rect 3148 5244 3200 5296
rect 3332 5244 3384 5296
rect 3424 5219 3476 5228
rect 3424 5185 3433 5219
rect 3433 5185 3467 5219
rect 3467 5185 3476 5219
rect 3424 5176 3476 5185
rect 4528 5287 4580 5296
rect 4528 5253 4537 5287
rect 4537 5253 4571 5287
rect 4571 5253 4580 5287
rect 4528 5244 4580 5253
rect 5264 5244 5316 5296
rect 7748 5312 7800 5364
rect 10140 5312 10192 5364
rect 1584 5151 1636 5160
rect 1584 5117 1593 5151
rect 1593 5117 1627 5151
rect 1627 5117 1636 5151
rect 1584 5108 1636 5117
rect 4160 5108 4212 5160
rect 5080 5108 5132 5160
rect 6552 5151 6604 5160
rect 6552 5117 6561 5151
rect 6561 5117 6595 5151
rect 6595 5117 6604 5151
rect 6552 5108 6604 5117
rect 12440 5312 12492 5364
rect 14004 5355 14056 5364
rect 14004 5321 14013 5355
rect 14013 5321 14047 5355
rect 14047 5321 14056 5355
rect 14004 5312 14056 5321
rect 15568 5312 15620 5364
rect 12532 5244 12584 5296
rect 11520 5219 11572 5228
rect 11520 5185 11529 5219
rect 11529 5185 11563 5219
rect 11563 5185 11572 5219
rect 11520 5176 11572 5185
rect 14096 5176 14148 5228
rect 14464 5244 14516 5296
rect 14648 5244 14700 5296
rect 16396 5176 16448 5228
rect 3332 5083 3384 5092
rect 3332 5049 3341 5083
rect 3341 5049 3375 5083
rect 3375 5049 3384 5083
rect 3332 5040 3384 5049
rect 7564 5108 7616 5160
rect 7288 5040 7340 5092
rect 8208 5108 8260 5160
rect 10600 5151 10652 5160
rect 10600 5117 10609 5151
rect 10609 5117 10643 5151
rect 10643 5117 10652 5151
rect 10600 5108 10652 5117
rect 14556 5151 14608 5160
rect 14556 5117 14565 5151
rect 14565 5117 14599 5151
rect 14599 5117 14608 5151
rect 14556 5108 14608 5117
rect 15752 5108 15804 5160
rect 6368 5015 6420 5024
rect 6368 4981 6377 5015
rect 6377 4981 6411 5015
rect 6411 4981 6420 5015
rect 6368 4972 6420 4981
rect 14280 4972 14332 5024
rect 2985 4870 3037 4922
rect 3049 4870 3101 4922
rect 3113 4870 3165 4922
rect 3177 4870 3229 4922
rect 3241 4870 3293 4922
rect 7056 4870 7108 4922
rect 7120 4870 7172 4922
rect 7184 4870 7236 4922
rect 7248 4870 7300 4922
rect 7312 4870 7364 4922
rect 11127 4870 11179 4922
rect 11191 4870 11243 4922
rect 11255 4870 11307 4922
rect 11319 4870 11371 4922
rect 11383 4870 11435 4922
rect 15198 4870 15250 4922
rect 15262 4870 15314 4922
rect 15326 4870 15378 4922
rect 15390 4870 15442 4922
rect 15454 4870 15506 4922
rect 6920 4768 6972 4820
rect 7564 4811 7616 4820
rect 7564 4777 7573 4811
rect 7573 4777 7607 4811
rect 7607 4777 7616 4811
rect 7564 4768 7616 4777
rect 14556 4811 14608 4820
rect 14556 4777 14565 4811
rect 14565 4777 14599 4811
rect 14599 4777 14608 4811
rect 14556 4768 14608 4777
rect 5080 4675 5132 4684
rect 5080 4641 5089 4675
rect 5089 4641 5123 4675
rect 5123 4641 5132 4675
rect 5080 4632 5132 4641
rect 6368 4632 6420 4684
rect 6552 4632 6604 4684
rect 7380 4632 7432 4684
rect 14096 4700 14148 4752
rect 14464 4700 14516 4752
rect 16764 4675 16816 4684
rect 16764 4641 16773 4675
rect 16773 4641 16807 4675
rect 16807 4641 16816 4675
rect 16764 4632 16816 4641
rect 14004 4564 14056 4616
rect 14280 4607 14332 4616
rect 14280 4573 14289 4607
rect 14289 4573 14323 4607
rect 14323 4573 14332 4607
rect 14280 4564 14332 4573
rect 5264 4428 5316 4480
rect 10232 4496 10284 4548
rect 15752 4496 15804 4548
rect 15292 4471 15344 4480
rect 15292 4437 15301 4471
rect 15301 4437 15335 4471
rect 15335 4437 15344 4471
rect 15292 4428 15344 4437
rect 3645 4326 3697 4378
rect 3709 4326 3761 4378
rect 3773 4326 3825 4378
rect 3837 4326 3889 4378
rect 3901 4326 3953 4378
rect 7716 4326 7768 4378
rect 7780 4326 7832 4378
rect 7844 4326 7896 4378
rect 7908 4326 7960 4378
rect 7972 4326 8024 4378
rect 11787 4326 11839 4378
rect 11851 4326 11903 4378
rect 11915 4326 11967 4378
rect 11979 4326 12031 4378
rect 12043 4326 12095 4378
rect 15858 4326 15910 4378
rect 15922 4326 15974 4378
rect 15986 4326 16038 4378
rect 16050 4326 16102 4378
rect 16114 4326 16166 4378
rect 5172 4224 5224 4276
rect 5816 4224 5868 4276
rect 7564 4156 7616 4208
rect 5080 4131 5132 4140
rect 5080 4097 5089 4131
rect 5089 4097 5123 4131
rect 5123 4097 5132 4131
rect 5080 4088 5132 4097
rect 5448 4088 5500 4140
rect 8208 4131 8260 4140
rect 8208 4097 8217 4131
rect 8217 4097 8251 4131
rect 8251 4097 8260 4131
rect 8208 4088 8260 4097
rect 10232 4199 10284 4208
rect 10232 4165 10241 4199
rect 10241 4165 10275 4199
rect 10275 4165 10284 4199
rect 10232 4156 10284 4165
rect 12992 4156 13044 4208
rect 12624 4088 12676 4140
rect 12716 4131 12768 4140
rect 12716 4097 12725 4131
rect 12725 4097 12759 4131
rect 12759 4097 12768 4131
rect 12716 4088 12768 4097
rect 13452 4088 13504 4140
rect 8944 4020 8996 4072
rect 10048 3952 10100 4004
rect 15292 4088 15344 4140
rect 15476 4131 15528 4140
rect 15476 4097 15485 4131
rect 15485 4097 15519 4131
rect 15519 4097 15528 4131
rect 15476 4088 15528 4097
rect 15568 4131 15620 4140
rect 15568 4097 15577 4131
rect 15577 4097 15611 4131
rect 15611 4097 15620 4131
rect 15568 4088 15620 4097
rect 16580 4088 16632 4140
rect 16488 3952 16540 4004
rect 4712 3884 4764 3936
rect 9864 3884 9916 3936
rect 12256 3884 12308 3936
rect 14096 3884 14148 3936
rect 15660 3884 15712 3936
rect 2985 3782 3037 3834
rect 3049 3782 3101 3834
rect 3113 3782 3165 3834
rect 3177 3782 3229 3834
rect 3241 3782 3293 3834
rect 7056 3782 7108 3834
rect 7120 3782 7172 3834
rect 7184 3782 7236 3834
rect 7248 3782 7300 3834
rect 7312 3782 7364 3834
rect 11127 3782 11179 3834
rect 11191 3782 11243 3834
rect 11255 3782 11307 3834
rect 11319 3782 11371 3834
rect 11383 3782 11435 3834
rect 15198 3782 15250 3834
rect 15262 3782 15314 3834
rect 15326 3782 15378 3834
rect 15390 3782 15442 3834
rect 15454 3782 15506 3834
rect 5080 3680 5132 3732
rect 4160 3544 4212 3596
rect 5264 3544 5316 3596
rect 8116 3680 8168 3732
rect 8944 3723 8996 3732
rect 8944 3689 8953 3723
rect 8953 3689 8987 3723
rect 8987 3689 8996 3723
rect 8944 3680 8996 3689
rect 12624 3723 12676 3732
rect 12624 3689 12633 3723
rect 12633 3689 12667 3723
rect 12667 3689 12676 3723
rect 12624 3680 12676 3689
rect 12900 3723 12952 3732
rect 12900 3689 12909 3723
rect 12909 3689 12943 3723
rect 12943 3689 12952 3723
rect 12900 3680 12952 3689
rect 8208 3544 8260 3596
rect 4068 3451 4120 3460
rect 4068 3417 4077 3451
rect 4077 3417 4111 3451
rect 4111 3417 4120 3451
rect 4068 3408 4120 3417
rect 5448 3408 5500 3460
rect 5816 3451 5868 3460
rect 5816 3417 5825 3451
rect 5825 3417 5859 3451
rect 5859 3417 5868 3451
rect 5816 3408 5868 3417
rect 6276 3451 6328 3460
rect 6276 3417 6285 3451
rect 6285 3417 6319 3451
rect 6319 3417 6328 3451
rect 6276 3408 6328 3417
rect 7564 3408 7616 3460
rect 9036 3476 9088 3528
rect 11520 3544 11572 3596
rect 9864 3519 9916 3528
rect 9864 3485 9873 3519
rect 9873 3485 9907 3519
rect 9907 3485 9916 3519
rect 9864 3476 9916 3485
rect 10048 3519 10100 3528
rect 10048 3485 10057 3519
rect 10057 3485 10091 3519
rect 10091 3485 10100 3519
rect 10048 3476 10100 3485
rect 10140 3519 10192 3528
rect 10140 3485 10149 3519
rect 10149 3485 10183 3519
rect 10183 3485 10192 3519
rect 10140 3476 10192 3485
rect 10692 3476 10744 3528
rect 13452 3519 13504 3528
rect 13452 3485 13461 3519
rect 13461 3485 13495 3519
rect 13495 3485 13504 3519
rect 13452 3476 13504 3485
rect 13728 3680 13780 3732
rect 16580 3723 16632 3732
rect 16580 3689 16589 3723
rect 16589 3689 16623 3723
rect 16623 3689 16632 3723
rect 16580 3680 16632 3689
rect 14464 3544 14516 3596
rect 11152 3451 11204 3460
rect 11152 3417 11161 3451
rect 11161 3417 11195 3451
rect 11195 3417 11204 3451
rect 11152 3408 11204 3417
rect 6092 3340 6144 3392
rect 8668 3383 8720 3392
rect 8668 3349 8677 3383
rect 8677 3349 8711 3383
rect 8711 3349 8720 3383
rect 8668 3340 8720 3349
rect 11612 3408 11664 3460
rect 12992 3408 13044 3460
rect 14648 3408 14700 3460
rect 12900 3340 12952 3392
rect 13360 3383 13412 3392
rect 13360 3349 13369 3383
rect 13369 3349 13403 3383
rect 13403 3349 13412 3383
rect 13360 3340 13412 3349
rect 13636 3340 13688 3392
rect 15384 3340 15436 3392
rect 15844 3408 15896 3460
rect 16304 3519 16356 3528
rect 16304 3485 16313 3519
rect 16313 3485 16347 3519
rect 16347 3485 16356 3519
rect 16304 3476 16356 3485
rect 16856 3612 16908 3664
rect 17040 3519 17092 3528
rect 17040 3485 17049 3519
rect 17049 3485 17083 3519
rect 17083 3485 17092 3519
rect 17040 3476 17092 3485
rect 15752 3340 15804 3392
rect 3645 3238 3697 3290
rect 3709 3238 3761 3290
rect 3773 3238 3825 3290
rect 3837 3238 3889 3290
rect 3901 3238 3953 3290
rect 7716 3238 7768 3290
rect 7780 3238 7832 3290
rect 7844 3238 7896 3290
rect 7908 3238 7960 3290
rect 7972 3238 8024 3290
rect 11787 3238 11839 3290
rect 11851 3238 11903 3290
rect 11915 3238 11967 3290
rect 11979 3238 12031 3290
rect 12043 3238 12095 3290
rect 15858 3238 15910 3290
rect 15922 3238 15974 3290
rect 15986 3238 16038 3290
rect 16050 3238 16102 3290
rect 16114 3238 16166 3290
rect 4068 3136 4120 3188
rect 4712 3136 4764 3188
rect 5724 3136 5776 3188
rect 6276 3136 6328 3188
rect 7564 3068 7616 3120
rect 9036 3179 9088 3188
rect 9036 3145 9045 3179
rect 9045 3145 9079 3179
rect 9079 3145 9088 3179
rect 9036 3136 9088 3145
rect 11152 3136 11204 3188
rect 4712 3043 4764 3052
rect 4712 3009 4721 3043
rect 4721 3009 4755 3043
rect 4755 3009 4764 3043
rect 4712 3000 4764 3009
rect 5356 2975 5408 2984
rect 5356 2941 5365 2975
rect 5365 2941 5399 2975
rect 5399 2941 5408 2975
rect 5356 2932 5408 2941
rect 5724 3000 5776 3052
rect 6092 3043 6144 3052
rect 6092 3009 6101 3043
rect 6101 3009 6135 3043
rect 6135 3009 6144 3043
rect 6092 3000 6144 3009
rect 8208 3000 8260 3052
rect 11612 3068 11664 3120
rect 13360 3136 13412 3188
rect 14648 3179 14700 3188
rect 14648 3145 14657 3179
rect 14657 3145 14691 3179
rect 14691 3145 14700 3179
rect 14648 3136 14700 3145
rect 16580 3136 16632 3188
rect 11520 3000 11572 3052
rect 12256 3043 12308 3052
rect 12256 3009 12265 3043
rect 12265 3009 12299 3043
rect 12299 3009 12308 3043
rect 12256 3000 12308 3009
rect 13636 3068 13688 3120
rect 14096 3111 14148 3120
rect 14096 3077 14105 3111
rect 14105 3077 14139 3111
rect 14139 3077 14148 3111
rect 14096 3068 14148 3077
rect 14464 3000 14516 3052
rect 15752 3068 15804 3120
rect 15200 3000 15252 3052
rect 15660 3043 15712 3052
rect 15660 3009 15669 3043
rect 15669 3009 15703 3043
rect 15703 3009 15712 3043
rect 15660 3000 15712 3009
rect 17040 3043 17092 3052
rect 17040 3009 17049 3043
rect 17049 3009 17083 3043
rect 17083 3009 17092 3043
rect 17040 3000 17092 3009
rect 8668 2975 8720 2984
rect 8668 2941 8677 2975
rect 8677 2941 8711 2975
rect 8711 2941 8720 2975
rect 8668 2932 8720 2941
rect 11888 2932 11940 2984
rect 11520 2864 11572 2916
rect 15384 2864 15436 2916
rect 15568 2864 15620 2916
rect 5356 2796 5408 2848
rect 11980 2796 12032 2848
rect 2985 2694 3037 2746
rect 3049 2694 3101 2746
rect 3113 2694 3165 2746
rect 3177 2694 3229 2746
rect 3241 2694 3293 2746
rect 7056 2694 7108 2746
rect 7120 2694 7172 2746
rect 7184 2694 7236 2746
rect 7248 2694 7300 2746
rect 7312 2694 7364 2746
rect 11127 2694 11179 2746
rect 11191 2694 11243 2746
rect 11255 2694 11307 2746
rect 11319 2694 11371 2746
rect 11383 2694 11435 2746
rect 15198 2694 15250 2746
rect 15262 2694 15314 2746
rect 15326 2694 15378 2746
rect 15390 2694 15442 2746
rect 15454 2694 15506 2746
rect 5448 2635 5500 2644
rect 5448 2601 5457 2635
rect 5457 2601 5491 2635
rect 5491 2601 5500 2635
rect 5448 2592 5500 2601
rect 6828 2592 6880 2644
rect 8300 2592 8352 2644
rect 10140 2592 10192 2644
rect 10232 2592 10284 2644
rect 11612 2592 11664 2644
rect 13452 2592 13504 2644
rect 11520 2567 11572 2576
rect 11520 2533 11529 2567
rect 11529 2533 11563 2567
rect 11563 2533 11572 2567
rect 11520 2524 11572 2533
rect 11980 2499 12032 2508
rect 11980 2465 11989 2499
rect 11989 2465 12023 2499
rect 12023 2465 12032 2499
rect 11980 2456 12032 2465
rect 5172 2388 5224 2440
rect 7104 2388 7156 2440
rect 8392 2388 8444 2440
rect 9680 2388 9732 2440
rect 10324 2388 10376 2440
rect 10968 2388 11020 2440
rect 11888 2431 11940 2440
rect 11888 2397 11897 2431
rect 11897 2397 11931 2431
rect 11931 2397 11940 2431
rect 11888 2388 11940 2397
rect 12900 2388 12952 2440
rect 3645 2150 3697 2202
rect 3709 2150 3761 2202
rect 3773 2150 3825 2202
rect 3837 2150 3889 2202
rect 3901 2150 3953 2202
rect 7716 2150 7768 2202
rect 7780 2150 7832 2202
rect 7844 2150 7896 2202
rect 7908 2150 7960 2202
rect 7972 2150 8024 2202
rect 11787 2150 11839 2202
rect 11851 2150 11903 2202
rect 11915 2150 11967 2202
rect 11979 2150 12031 2202
rect 12043 2150 12095 2202
rect 15858 2150 15910 2202
rect 15922 2150 15974 2202
rect 15986 2150 16038 2202
rect 16050 2150 16102 2202
rect 16114 2150 16166 2202
<< metal2 >>
rect 5170 19860 5226 20660
rect 8390 19860 8446 20660
rect 9034 19860 9090 20660
rect 9678 19860 9734 20660
rect 10966 19860 11022 20660
rect 12254 19860 12310 20660
rect 2985 17980 3293 17989
rect 2985 17978 2991 17980
rect 3047 17978 3071 17980
rect 3127 17978 3151 17980
rect 3207 17978 3231 17980
rect 3287 17978 3293 17980
rect 3047 17926 3049 17978
rect 3229 17926 3231 17978
rect 2985 17924 2991 17926
rect 3047 17924 3071 17926
rect 3127 17924 3151 17926
rect 3207 17924 3231 17926
rect 3287 17924 3293 17926
rect 2985 17915 3293 17924
rect 5080 17808 5132 17814
rect 5080 17750 5132 17756
rect 4068 17672 4120 17678
rect 4068 17614 4120 17620
rect 3645 17436 3953 17445
rect 3645 17434 3651 17436
rect 3707 17434 3731 17436
rect 3787 17434 3811 17436
rect 3867 17434 3891 17436
rect 3947 17434 3953 17436
rect 3707 17382 3709 17434
rect 3889 17382 3891 17434
rect 3645 17380 3651 17382
rect 3707 17380 3731 17382
rect 3787 17380 3811 17382
rect 3867 17380 3891 17382
rect 3947 17380 3953 17382
rect 3645 17371 3953 17380
rect 846 17232 902 17241
rect 846 17167 848 17176
rect 900 17167 902 17176
rect 848 17138 900 17144
rect 3424 17128 3476 17134
rect 3424 17070 3476 17076
rect 1584 16992 1636 16998
rect 1584 16934 1636 16940
rect 1596 16590 1624 16934
rect 2985 16892 3293 16901
rect 2985 16890 2991 16892
rect 3047 16890 3071 16892
rect 3127 16890 3151 16892
rect 3207 16890 3231 16892
rect 3287 16890 3293 16892
rect 3047 16838 3049 16890
rect 3229 16838 3231 16890
rect 2985 16836 2991 16838
rect 3047 16836 3071 16838
rect 3127 16836 3151 16838
rect 3207 16836 3231 16838
rect 3287 16836 3293 16838
rect 2985 16827 3293 16836
rect 1584 16584 1636 16590
rect 1584 16526 1636 16532
rect 1584 16448 1636 16454
rect 1584 16390 1636 16396
rect 1400 16040 1452 16046
rect 1400 15982 1452 15988
rect 1030 15736 1086 15745
rect 1030 15671 1086 15680
rect 1044 15502 1072 15671
rect 1412 15638 1440 15982
rect 1400 15632 1452 15638
rect 1400 15574 1452 15580
rect 1032 15496 1084 15502
rect 1032 15438 1084 15444
rect 1412 14634 1440 15574
rect 1596 15434 1624 16390
rect 3332 16108 3384 16114
rect 3332 16050 3384 16056
rect 1676 16040 1728 16046
rect 1676 15982 1728 15988
rect 1688 15706 1716 15982
rect 2780 15904 2832 15910
rect 2780 15846 2832 15852
rect 1676 15700 1728 15706
rect 1676 15642 1728 15648
rect 2792 15450 2820 15846
rect 2985 15804 3293 15813
rect 2985 15802 2991 15804
rect 3047 15802 3071 15804
rect 3127 15802 3151 15804
rect 3207 15802 3231 15804
rect 3287 15802 3293 15804
rect 3047 15750 3049 15802
rect 3229 15750 3231 15802
rect 2985 15748 2991 15750
rect 3047 15748 3071 15750
rect 3127 15748 3151 15750
rect 3207 15748 3231 15750
rect 3287 15748 3293 15750
rect 2985 15739 3293 15748
rect 3240 15700 3292 15706
rect 3240 15642 3292 15648
rect 3252 15570 3280 15642
rect 3240 15564 3292 15570
rect 3240 15506 3292 15512
rect 2700 15434 2820 15450
rect 2872 15496 2924 15502
rect 2872 15438 2924 15444
rect 2964 15496 3016 15502
rect 2964 15438 3016 15444
rect 1584 15428 1636 15434
rect 1584 15370 1636 15376
rect 2688 15428 2820 15434
rect 2740 15422 2820 15428
rect 2688 15370 2740 15376
rect 1412 14606 1532 14634
rect 1400 13932 1452 13938
rect 1400 13874 1452 13880
rect 1412 13705 1440 13874
rect 1398 13696 1454 13705
rect 1398 13631 1454 13640
rect 1504 13546 1532 14606
rect 1412 13518 1532 13546
rect 848 13320 900 13326
rect 848 13262 900 13268
rect 860 13161 888 13262
rect 846 13152 902 13161
rect 846 13087 902 13096
rect 1412 12850 1440 13518
rect 1400 12844 1452 12850
rect 1400 12786 1452 12792
rect 1412 11218 1440 12786
rect 1400 11212 1452 11218
rect 1400 11154 1452 11160
rect 1412 11014 1440 11154
rect 1400 11008 1452 11014
rect 1400 10950 1452 10956
rect 846 10840 902 10849
rect 846 10775 902 10784
rect 860 10674 888 10775
rect 848 10668 900 10674
rect 848 10610 900 10616
rect 1400 10056 1452 10062
rect 1400 9998 1452 10004
rect 1412 9625 1440 9998
rect 1596 9654 1624 15370
rect 2792 15094 2820 15422
rect 2780 15088 2832 15094
rect 2780 15030 2832 15036
rect 2884 15026 2912 15438
rect 2976 15162 3004 15438
rect 3252 15178 3280 15506
rect 3344 15366 3372 16050
rect 3436 15638 3464 17070
rect 3645 16348 3953 16357
rect 3645 16346 3651 16348
rect 3707 16346 3731 16348
rect 3787 16346 3811 16348
rect 3867 16346 3891 16348
rect 3947 16346 3953 16348
rect 3707 16294 3709 16346
rect 3889 16294 3891 16346
rect 3645 16292 3651 16294
rect 3707 16292 3731 16294
rect 3787 16292 3811 16294
rect 3867 16292 3891 16294
rect 3947 16292 3953 16294
rect 3645 16283 3953 16292
rect 3516 16108 3568 16114
rect 3516 16050 3568 16056
rect 3424 15632 3476 15638
rect 3424 15574 3476 15580
rect 3332 15360 3384 15366
rect 3332 15302 3384 15308
rect 2964 15156 3016 15162
rect 3252 15150 3372 15178
rect 3528 15162 3556 16050
rect 3884 15904 3936 15910
rect 3884 15846 3936 15852
rect 3896 15570 3924 15846
rect 4080 15706 4108 17614
rect 5092 17610 5120 17750
rect 5184 17746 5212 19860
rect 7056 17980 7364 17989
rect 7056 17978 7062 17980
rect 7118 17978 7142 17980
rect 7198 17978 7222 17980
rect 7278 17978 7302 17980
rect 7358 17978 7364 17980
rect 7118 17926 7120 17978
rect 7300 17926 7302 17978
rect 7056 17924 7062 17926
rect 7118 17924 7142 17926
rect 7198 17924 7222 17926
rect 7278 17924 7302 17926
rect 7358 17924 7364 17926
rect 7056 17915 7364 17924
rect 5172 17740 5224 17746
rect 5172 17682 5224 17688
rect 8404 17678 8432 19860
rect 8944 17808 8996 17814
rect 8944 17750 8996 17756
rect 8956 17678 8984 17750
rect 9048 17746 9076 19860
rect 9588 17876 9640 17882
rect 9588 17818 9640 17824
rect 9036 17740 9088 17746
rect 9036 17682 9088 17688
rect 9404 17740 9456 17746
rect 9404 17682 9456 17688
rect 5448 17672 5500 17678
rect 5448 17614 5500 17620
rect 8392 17672 8444 17678
rect 8392 17614 8444 17620
rect 8944 17672 8996 17678
rect 8944 17614 8996 17620
rect 9128 17672 9180 17678
rect 9128 17614 9180 17620
rect 5080 17604 5132 17610
rect 5080 17546 5132 17552
rect 5264 17604 5316 17610
rect 5264 17546 5316 17552
rect 4160 17264 4212 17270
rect 4160 17206 4212 17212
rect 4172 16182 4200 17206
rect 5092 16590 5120 17546
rect 5276 16998 5304 17546
rect 5460 17202 5488 17614
rect 5908 17604 5960 17610
rect 5908 17546 5960 17552
rect 5540 17536 5592 17542
rect 5540 17478 5592 17484
rect 5552 17270 5580 17478
rect 5920 17338 5948 17546
rect 8484 17536 8536 17542
rect 8484 17478 8536 17484
rect 8576 17536 8628 17542
rect 8576 17478 8628 17484
rect 8668 17536 8720 17542
rect 8668 17478 8720 17484
rect 8956 17490 8984 17614
rect 7716 17436 8024 17445
rect 7716 17434 7722 17436
rect 7778 17434 7802 17436
rect 7858 17434 7882 17436
rect 7938 17434 7962 17436
rect 8018 17434 8024 17436
rect 7778 17382 7780 17434
rect 7960 17382 7962 17434
rect 7716 17380 7722 17382
rect 7778 17380 7802 17382
rect 7858 17380 7882 17382
rect 7938 17380 7962 17382
rect 8018 17380 8024 17382
rect 7716 17371 8024 17380
rect 5908 17332 5960 17338
rect 5908 17274 5960 17280
rect 5540 17264 5592 17270
rect 5540 17206 5592 17212
rect 5448 17196 5500 17202
rect 5448 17138 5500 17144
rect 6000 17196 6052 17202
rect 6000 17138 6052 17144
rect 6736 17196 6788 17202
rect 6736 17138 6788 17144
rect 8392 17196 8444 17202
rect 8392 17138 8444 17144
rect 5264 16992 5316 16998
rect 5264 16934 5316 16940
rect 5276 16590 5304 16934
rect 5460 16794 5488 17138
rect 6012 16794 6040 17138
rect 6276 17128 6328 17134
rect 6276 17070 6328 17076
rect 6552 17128 6604 17134
rect 6748 17082 6776 17138
rect 6604 17076 6776 17082
rect 6552 17070 6776 17076
rect 6092 16992 6144 16998
rect 6092 16934 6144 16940
rect 5448 16788 5500 16794
rect 5448 16730 5500 16736
rect 6000 16788 6052 16794
rect 6000 16730 6052 16736
rect 5080 16584 5132 16590
rect 5080 16526 5132 16532
rect 5264 16584 5316 16590
rect 5264 16526 5316 16532
rect 6012 16522 6040 16730
rect 6104 16658 6132 16934
rect 6092 16652 6144 16658
rect 6092 16594 6144 16600
rect 6000 16516 6052 16522
rect 6000 16458 6052 16464
rect 5080 16448 5132 16454
rect 5080 16390 5132 16396
rect 4160 16176 4212 16182
rect 4160 16118 4212 16124
rect 4068 15700 4120 15706
rect 4068 15642 4120 15648
rect 3884 15564 3936 15570
rect 3884 15506 3936 15512
rect 3976 15496 4028 15502
rect 3976 15438 4028 15444
rect 3645 15260 3953 15269
rect 3645 15258 3651 15260
rect 3707 15258 3731 15260
rect 3787 15258 3811 15260
rect 3867 15258 3891 15260
rect 3947 15258 3953 15260
rect 3707 15206 3709 15258
rect 3889 15206 3891 15258
rect 3645 15204 3651 15206
rect 3707 15204 3731 15206
rect 3787 15204 3811 15206
rect 3867 15204 3891 15206
rect 3947 15204 3953 15206
rect 3645 15195 3953 15204
rect 2964 15098 3016 15104
rect 2872 15020 2924 15026
rect 2872 14962 2924 14968
rect 2985 14716 3293 14725
rect 2985 14714 2991 14716
rect 3047 14714 3071 14716
rect 3127 14714 3151 14716
rect 3207 14714 3231 14716
rect 3287 14714 3293 14716
rect 3047 14662 3049 14714
rect 3229 14662 3231 14714
rect 2985 14660 2991 14662
rect 3047 14660 3071 14662
rect 3127 14660 3151 14662
rect 3207 14660 3231 14662
rect 3287 14660 3293 14662
rect 2985 14651 3293 14660
rect 2780 14068 2832 14074
rect 2780 14010 2832 14016
rect 2792 13394 2820 14010
rect 2985 13628 3293 13637
rect 2985 13626 2991 13628
rect 3047 13626 3071 13628
rect 3127 13626 3151 13628
rect 3207 13626 3231 13628
rect 3287 13626 3293 13628
rect 3047 13574 3049 13626
rect 3229 13574 3231 13626
rect 2985 13572 2991 13574
rect 3047 13572 3071 13574
rect 3127 13572 3151 13574
rect 3207 13572 3231 13574
rect 3287 13572 3293 13574
rect 2985 13563 3293 13572
rect 3344 13394 3372 15150
rect 3516 15156 3568 15162
rect 3516 15098 3568 15104
rect 3516 14952 3568 14958
rect 3516 14894 3568 14900
rect 2780 13388 2832 13394
rect 2780 13330 2832 13336
rect 3332 13388 3384 13394
rect 3332 13330 3384 13336
rect 3240 13252 3292 13258
rect 3240 13194 3292 13200
rect 2688 13184 2740 13190
rect 2688 13126 2740 13132
rect 1676 12776 1728 12782
rect 1676 12718 1728 12724
rect 1688 12442 1716 12718
rect 1676 12436 1728 12442
rect 1676 12378 1728 12384
rect 2700 12238 2728 13126
rect 3252 12986 3280 13194
rect 3528 13190 3556 14894
rect 3988 14618 4016 15438
rect 5092 14958 5120 16390
rect 5172 16176 5224 16182
rect 5172 16118 5224 16124
rect 5184 15434 5212 16118
rect 5264 15564 5316 15570
rect 5264 15506 5316 15512
rect 5172 15428 5224 15434
rect 5172 15370 5224 15376
rect 5080 14952 5132 14958
rect 5080 14894 5132 14900
rect 3976 14612 4028 14618
rect 3976 14554 4028 14560
rect 5184 14346 5212 15370
rect 5276 14482 5304 15506
rect 6104 15026 6132 16594
rect 6288 15706 6316 17070
rect 6564 17054 6776 17070
rect 6460 16992 6512 16998
rect 6460 16934 6512 16940
rect 6472 16658 6500 16934
rect 7056 16892 7364 16901
rect 7056 16890 7062 16892
rect 7118 16890 7142 16892
rect 7198 16890 7222 16892
rect 7278 16890 7302 16892
rect 7358 16890 7364 16892
rect 7118 16838 7120 16890
rect 7300 16838 7302 16890
rect 7056 16836 7062 16838
rect 7118 16836 7142 16838
rect 7198 16836 7222 16838
rect 7278 16836 7302 16838
rect 7358 16836 7364 16838
rect 7056 16827 7364 16836
rect 6460 16652 6512 16658
rect 6460 16594 6512 16600
rect 8404 16590 8432 17138
rect 8392 16584 8444 16590
rect 8392 16526 8444 16532
rect 8208 16516 8260 16522
rect 8208 16458 8260 16464
rect 8116 16448 8168 16454
rect 8116 16390 8168 16396
rect 7716 16348 8024 16357
rect 7716 16346 7722 16348
rect 7778 16346 7802 16348
rect 7858 16346 7882 16348
rect 7938 16346 7962 16348
rect 8018 16346 8024 16348
rect 7778 16294 7780 16346
rect 7960 16294 7962 16346
rect 7716 16292 7722 16294
rect 7778 16292 7802 16294
rect 7858 16292 7882 16294
rect 7938 16292 7962 16294
rect 8018 16292 8024 16294
rect 7716 16283 8024 16292
rect 7056 15804 7364 15813
rect 7056 15802 7062 15804
rect 7118 15802 7142 15804
rect 7198 15802 7222 15804
rect 7278 15802 7302 15804
rect 7358 15802 7364 15804
rect 7118 15750 7120 15802
rect 7300 15750 7302 15802
rect 7056 15748 7062 15750
rect 7118 15748 7142 15750
rect 7198 15748 7222 15750
rect 7278 15748 7302 15750
rect 7358 15748 7364 15750
rect 7056 15739 7364 15748
rect 6276 15700 6328 15706
rect 6276 15642 6328 15648
rect 7564 15496 7616 15502
rect 7564 15438 7616 15444
rect 7472 15428 7524 15434
rect 7472 15370 7524 15376
rect 7012 15360 7064 15366
rect 7012 15302 7064 15308
rect 7024 15094 7052 15302
rect 7012 15088 7064 15094
rect 7012 15030 7064 15036
rect 6092 15020 6144 15026
rect 6092 14962 6144 14968
rect 6104 14498 6132 14962
rect 7484 14958 7512 15370
rect 7472 14952 7524 14958
rect 7472 14894 7524 14900
rect 7380 14816 7432 14822
rect 7380 14758 7432 14764
rect 7056 14716 7364 14725
rect 7056 14714 7062 14716
rect 7118 14714 7142 14716
rect 7198 14714 7222 14716
rect 7278 14714 7302 14716
rect 7358 14714 7364 14716
rect 7118 14662 7120 14714
rect 7300 14662 7302 14714
rect 7056 14660 7062 14662
rect 7118 14660 7142 14662
rect 7198 14660 7222 14662
rect 7278 14660 7302 14662
rect 7358 14660 7364 14662
rect 7056 14651 7364 14660
rect 7392 14550 7420 14758
rect 7484 14618 7512 14894
rect 7576 14822 7604 15438
rect 7716 15260 8024 15269
rect 7716 15258 7722 15260
rect 7778 15258 7802 15260
rect 7858 15258 7882 15260
rect 7938 15258 7962 15260
rect 8018 15258 8024 15260
rect 7778 15206 7780 15258
rect 7960 15206 7962 15258
rect 7716 15204 7722 15206
rect 7778 15204 7802 15206
rect 7858 15204 7882 15206
rect 7938 15204 7962 15206
rect 8018 15204 8024 15206
rect 7716 15195 8024 15204
rect 8128 15178 8156 16390
rect 8220 15570 8248 16458
rect 8208 15564 8260 15570
rect 8208 15506 8260 15512
rect 8300 15428 8352 15434
rect 8300 15370 8352 15376
rect 8128 15150 8248 15178
rect 8312 15162 8340 15370
rect 7564 14816 7616 14822
rect 7564 14758 7616 14764
rect 7472 14612 7524 14618
rect 7472 14554 7524 14560
rect 7380 14544 7432 14550
rect 6104 14482 6224 14498
rect 7380 14486 7432 14492
rect 7576 14482 7604 14758
rect 5264 14476 5316 14482
rect 5264 14418 5316 14424
rect 6092 14476 6224 14482
rect 6144 14470 6224 14476
rect 6092 14418 6144 14424
rect 5172 14340 5224 14346
rect 5172 14282 5224 14288
rect 3645 14172 3953 14181
rect 3645 14170 3651 14172
rect 3707 14170 3731 14172
rect 3787 14170 3811 14172
rect 3867 14170 3891 14172
rect 3947 14170 3953 14172
rect 3707 14118 3709 14170
rect 3889 14118 3891 14170
rect 3645 14116 3651 14118
rect 3707 14116 3731 14118
rect 3787 14116 3811 14118
rect 3867 14116 3891 14118
rect 3947 14116 3953 14118
rect 3645 14107 3953 14116
rect 3976 13320 4028 13326
rect 3976 13262 4028 13268
rect 3424 13184 3476 13190
rect 3424 13126 3476 13132
rect 3516 13184 3568 13190
rect 3516 13126 3568 13132
rect 3240 12980 3292 12986
rect 3240 12922 3292 12928
rect 2780 12844 2832 12850
rect 2780 12786 2832 12792
rect 2688 12232 2740 12238
rect 2688 12174 2740 12180
rect 2792 11150 2820 12786
rect 2872 12776 2924 12782
rect 2872 12718 2924 12724
rect 3332 12776 3384 12782
rect 3332 12718 3384 12724
rect 2884 12170 2912 12718
rect 2985 12540 3293 12549
rect 2985 12538 2991 12540
rect 3047 12538 3071 12540
rect 3127 12538 3151 12540
rect 3207 12538 3231 12540
rect 3287 12538 3293 12540
rect 3047 12486 3049 12538
rect 3229 12486 3231 12538
rect 2985 12484 2991 12486
rect 3047 12484 3071 12486
rect 3127 12484 3151 12486
rect 3207 12484 3231 12486
rect 3287 12484 3293 12486
rect 2985 12475 3293 12484
rect 3344 12442 3372 12718
rect 3332 12436 3384 12442
rect 3332 12378 3384 12384
rect 3436 12238 3464 13126
rect 3424 12232 3476 12238
rect 3424 12174 3476 12180
rect 2872 12164 2924 12170
rect 2872 12106 2924 12112
rect 2884 11354 2912 12106
rect 2985 11452 3293 11461
rect 2985 11450 2991 11452
rect 3047 11450 3071 11452
rect 3127 11450 3151 11452
rect 3207 11450 3231 11452
rect 3287 11450 3293 11452
rect 3047 11398 3049 11450
rect 3229 11398 3231 11450
rect 2985 11396 2991 11398
rect 3047 11396 3071 11398
rect 3127 11396 3151 11398
rect 3207 11396 3231 11398
rect 3287 11396 3293 11398
rect 2985 11387 3293 11396
rect 2872 11348 2924 11354
rect 2872 11290 2924 11296
rect 2780 11144 2832 11150
rect 2780 11086 2832 11092
rect 2596 11008 2648 11014
rect 2596 10950 2648 10956
rect 2608 10674 2636 10950
rect 2792 10810 2820 11086
rect 2780 10804 2832 10810
rect 2780 10746 2832 10752
rect 2044 10668 2096 10674
rect 2044 10610 2096 10616
rect 2596 10668 2648 10674
rect 2596 10610 2648 10616
rect 1584 9648 1636 9654
rect 1398 9616 1454 9625
rect 1584 9590 1636 9596
rect 1398 9551 1454 9560
rect 1596 9450 1624 9590
rect 2056 9518 2084 10610
rect 2872 10464 2924 10470
rect 2872 10406 2924 10412
rect 2884 9722 2912 10406
rect 2985 10364 3293 10373
rect 2985 10362 2991 10364
rect 3047 10362 3071 10364
rect 3127 10362 3151 10364
rect 3207 10362 3231 10364
rect 3287 10362 3293 10364
rect 3047 10310 3049 10362
rect 3229 10310 3231 10362
rect 2985 10308 2991 10310
rect 3047 10308 3071 10310
rect 3127 10308 3151 10310
rect 3207 10308 3231 10310
rect 3287 10308 3293 10310
rect 2985 10299 3293 10308
rect 2964 9920 3016 9926
rect 2964 9862 3016 9868
rect 2872 9716 2924 9722
rect 2872 9658 2924 9664
rect 2976 9625 3004 9862
rect 3528 9738 3556 13126
rect 3645 13084 3953 13093
rect 3645 13082 3651 13084
rect 3707 13082 3731 13084
rect 3787 13082 3811 13084
rect 3867 13082 3891 13084
rect 3947 13082 3953 13084
rect 3707 13030 3709 13082
rect 3889 13030 3891 13082
rect 3645 13028 3651 13030
rect 3707 13028 3731 13030
rect 3787 13028 3811 13030
rect 3867 13028 3891 13030
rect 3947 13028 3953 13030
rect 3645 13019 3953 13028
rect 3645 11996 3953 12005
rect 3645 11994 3651 11996
rect 3707 11994 3731 11996
rect 3787 11994 3811 11996
rect 3867 11994 3891 11996
rect 3947 11994 3953 11996
rect 3707 11942 3709 11994
rect 3889 11942 3891 11994
rect 3645 11940 3651 11942
rect 3707 11940 3731 11942
rect 3787 11940 3811 11942
rect 3867 11940 3891 11942
rect 3947 11940 3953 11942
rect 3645 11931 3953 11940
rect 3645 10908 3953 10917
rect 3645 10906 3651 10908
rect 3707 10906 3731 10908
rect 3787 10906 3811 10908
rect 3867 10906 3891 10908
rect 3947 10906 3953 10908
rect 3707 10854 3709 10906
rect 3889 10854 3891 10906
rect 3645 10852 3651 10854
rect 3707 10852 3731 10854
rect 3787 10852 3811 10854
rect 3867 10852 3891 10854
rect 3947 10852 3953 10854
rect 3645 10843 3953 10852
rect 3645 9820 3953 9829
rect 3645 9818 3651 9820
rect 3707 9818 3731 9820
rect 3787 9818 3811 9820
rect 3867 9818 3891 9820
rect 3947 9818 3953 9820
rect 3707 9766 3709 9818
rect 3889 9766 3891 9818
rect 3645 9764 3651 9766
rect 3707 9764 3731 9766
rect 3787 9764 3811 9766
rect 3867 9764 3891 9766
rect 3947 9764 3953 9766
rect 3645 9755 3953 9764
rect 3160 9710 3556 9738
rect 2962 9616 3018 9625
rect 2688 9580 2740 9586
rect 2688 9522 2740 9528
rect 2872 9580 2924 9586
rect 2962 9551 2964 9560
rect 2872 9522 2924 9528
rect 3016 9551 3018 9560
rect 2964 9522 3016 9528
rect 2044 9512 2096 9518
rect 2412 9512 2464 9518
rect 2044 9454 2096 9460
rect 2410 9480 2412 9489
rect 2464 9480 2466 9489
rect 1584 9444 1636 9450
rect 1584 9386 1636 9392
rect 1492 9376 1544 9382
rect 1492 9318 1544 9324
rect 1676 9376 1728 9382
rect 1676 9318 1728 9324
rect 1504 9194 1532 9318
rect 1504 9166 1624 9194
rect 1596 8838 1624 9166
rect 1688 9042 1716 9318
rect 1676 9036 1728 9042
rect 1676 8978 1728 8984
rect 1584 8832 1636 8838
rect 846 8800 902 8809
rect 1584 8774 1636 8780
rect 846 8735 902 8744
rect 860 8498 888 8735
rect 848 8492 900 8498
rect 848 8434 900 8440
rect 848 7880 900 7886
rect 848 7822 900 7828
rect 860 7721 888 7822
rect 846 7712 902 7721
rect 846 7647 902 7656
rect 1596 6730 1624 8774
rect 2056 8634 2084 9454
rect 2410 9415 2466 9424
rect 2700 9178 2728 9522
rect 2884 9466 2912 9522
rect 3160 9466 3188 9710
rect 3988 9654 4016 13262
rect 4712 13252 4764 13258
rect 4712 13194 4764 13200
rect 4724 12918 4752 13194
rect 5184 12918 5212 14282
rect 4712 12912 4764 12918
rect 4712 12854 4764 12860
rect 5172 12912 5224 12918
rect 5172 12854 5224 12860
rect 4436 12776 4488 12782
rect 4436 12718 4488 12724
rect 4068 12708 4120 12714
rect 4068 12650 4120 12656
rect 4080 12306 4108 12650
rect 4448 12434 4476 12718
rect 4356 12406 4476 12434
rect 4068 12300 4120 12306
rect 4068 12242 4120 12248
rect 4356 12170 4384 12406
rect 5184 12238 5212 12854
rect 5276 12782 5304 14418
rect 6092 14340 6144 14346
rect 6092 14282 6144 14288
rect 6104 14074 6132 14282
rect 6092 14068 6144 14074
rect 6092 14010 6144 14016
rect 5540 13932 5592 13938
rect 5540 13874 5592 13880
rect 5356 13864 5408 13870
rect 5356 13806 5408 13812
rect 5368 13530 5396 13806
rect 5356 13524 5408 13530
rect 5356 13466 5408 13472
rect 5552 13326 5580 13874
rect 5540 13320 5592 13326
rect 5540 13262 5592 13268
rect 5264 12776 5316 12782
rect 5264 12718 5316 12724
rect 5552 12442 5580 13262
rect 6196 12782 6224 14470
rect 7564 14476 7616 14482
rect 7564 14418 7616 14424
rect 7564 14340 7616 14346
rect 7564 14282 7616 14288
rect 7576 14074 7604 14282
rect 7716 14172 8024 14181
rect 7716 14170 7722 14172
rect 7778 14170 7802 14172
rect 7858 14170 7882 14172
rect 7938 14170 7962 14172
rect 8018 14170 8024 14172
rect 7778 14118 7780 14170
rect 7960 14118 7962 14170
rect 7716 14116 7722 14118
rect 7778 14116 7802 14118
rect 7858 14116 7882 14118
rect 7938 14116 7962 14118
rect 8018 14116 8024 14118
rect 7716 14107 8024 14116
rect 7564 14068 7616 14074
rect 7564 14010 7616 14016
rect 7056 13628 7364 13637
rect 7056 13626 7062 13628
rect 7118 13626 7142 13628
rect 7198 13626 7222 13628
rect 7278 13626 7302 13628
rect 7358 13626 7364 13628
rect 7118 13574 7120 13626
rect 7300 13574 7302 13626
rect 7056 13572 7062 13574
rect 7118 13572 7142 13574
rect 7198 13572 7222 13574
rect 7278 13572 7302 13574
rect 7358 13572 7364 13574
rect 7056 13563 7364 13572
rect 8116 13388 8168 13394
rect 8116 13330 8168 13336
rect 6276 13320 6328 13326
rect 6276 13262 6328 13268
rect 6368 13320 6420 13326
rect 6368 13262 6420 13268
rect 6920 13320 6972 13326
rect 6920 13262 6972 13268
rect 7380 13320 7432 13326
rect 7380 13262 7432 13268
rect 6288 12986 6316 13262
rect 6380 13190 6408 13262
rect 6368 13184 6420 13190
rect 6368 13126 6420 13132
rect 6460 13184 6512 13190
rect 6460 13126 6512 13132
rect 6276 12980 6328 12986
rect 6276 12922 6328 12928
rect 6184 12776 6236 12782
rect 6184 12718 6236 12724
rect 5540 12436 5592 12442
rect 5540 12378 5592 12384
rect 5172 12232 5224 12238
rect 5172 12174 5224 12180
rect 4344 12164 4396 12170
rect 4344 12106 4396 12112
rect 4252 11552 4304 11558
rect 4252 11494 4304 11500
rect 4264 11218 4292 11494
rect 4356 11218 4384 12106
rect 4712 11756 4764 11762
rect 4712 11698 4764 11704
rect 4252 11212 4304 11218
rect 4252 11154 4304 11160
rect 4344 11212 4396 11218
rect 4344 11154 4396 11160
rect 4160 11144 4212 11150
rect 4160 11086 4212 11092
rect 4172 10810 4200 11086
rect 4160 10804 4212 10810
rect 4160 10746 4212 10752
rect 4724 10606 4752 11698
rect 5184 11218 5212 12174
rect 6472 11898 6500 13126
rect 6828 12776 6880 12782
rect 6828 12718 6880 12724
rect 6000 11892 6052 11898
rect 6000 11834 6052 11840
rect 6460 11892 6512 11898
rect 6460 11834 6512 11840
rect 5816 11756 5868 11762
rect 5816 11698 5868 11704
rect 5908 11756 5960 11762
rect 5908 11698 5960 11704
rect 5356 11688 5408 11694
rect 5356 11630 5408 11636
rect 5172 11212 5224 11218
rect 5172 11154 5224 11160
rect 4804 11076 4856 11082
rect 4804 11018 4856 11024
rect 4816 10810 4844 11018
rect 5368 10810 5396 11630
rect 5828 11354 5856 11698
rect 5816 11348 5868 11354
rect 5816 11290 5868 11296
rect 4804 10804 4856 10810
rect 4804 10746 4856 10752
rect 5356 10804 5408 10810
rect 5356 10746 5408 10752
rect 5828 10674 5856 11290
rect 5816 10668 5868 10674
rect 5816 10610 5868 10616
rect 4712 10600 4764 10606
rect 4712 10542 4764 10548
rect 5920 10538 5948 11698
rect 5908 10532 5960 10538
rect 5908 10474 5960 10480
rect 3516 9648 3568 9654
rect 3422 9616 3478 9625
rect 3332 9580 3384 9586
rect 3516 9590 3568 9596
rect 3976 9648 4028 9654
rect 3976 9590 4028 9596
rect 3422 9551 3478 9560
rect 3332 9522 3384 9528
rect 3344 9489 3372 9522
rect 2792 9438 3188 9466
rect 3330 9480 3386 9489
rect 2688 9172 2740 9178
rect 2688 9114 2740 9120
rect 2044 8628 2096 8634
rect 2044 8570 2096 8576
rect 1676 8492 1728 8498
rect 1676 8434 1728 8440
rect 1688 8265 1716 8434
rect 2412 8288 2464 8294
rect 1674 8256 1730 8265
rect 2412 8230 2464 8236
rect 1674 8191 1730 8200
rect 2228 8084 2280 8090
rect 2228 8026 2280 8032
rect 2240 7410 2268 8026
rect 2424 7410 2452 8230
rect 2228 7404 2280 7410
rect 2228 7346 2280 7352
rect 2412 7404 2464 7410
rect 2412 7346 2464 7352
rect 1584 6724 1636 6730
rect 1584 6666 1636 6672
rect 1400 5704 1452 5710
rect 1400 5646 1452 5652
rect 1412 5545 1440 5646
rect 1398 5536 1454 5545
rect 1398 5471 1454 5480
rect 1596 5166 1624 6666
rect 2424 5710 2452 7346
rect 2792 6458 2820 9438
rect 3330 9415 3386 9424
rect 2985 9276 3293 9285
rect 2985 9274 2991 9276
rect 3047 9274 3071 9276
rect 3127 9274 3151 9276
rect 3207 9274 3231 9276
rect 3287 9274 3293 9276
rect 3047 9222 3049 9274
rect 3229 9222 3231 9274
rect 2985 9220 2991 9222
rect 3047 9220 3071 9222
rect 3127 9220 3151 9222
rect 3207 9220 3231 9222
rect 3287 9220 3293 9222
rect 2985 9211 3293 9220
rect 3344 9178 3372 9415
rect 3332 9172 3384 9178
rect 3332 9114 3384 9120
rect 3436 8974 3464 9551
rect 3528 8974 3556 9590
rect 5724 9580 5776 9586
rect 5724 9522 5776 9528
rect 5816 9580 5868 9586
rect 6012 9568 6040 11834
rect 6736 11756 6788 11762
rect 6736 11698 6788 11704
rect 6748 10810 6776 11698
rect 6840 11150 6868 12718
rect 6932 11762 6960 13262
rect 7056 12540 7364 12549
rect 7056 12538 7062 12540
rect 7118 12538 7142 12540
rect 7198 12538 7222 12540
rect 7278 12538 7302 12540
rect 7358 12538 7364 12540
rect 7118 12486 7120 12538
rect 7300 12486 7302 12538
rect 7056 12484 7062 12486
rect 7118 12484 7142 12486
rect 7198 12484 7222 12486
rect 7278 12484 7302 12486
rect 7358 12484 7364 12486
rect 7056 12475 7364 12484
rect 7392 12306 7420 13262
rect 7564 13184 7616 13190
rect 7564 13126 7616 13132
rect 7472 12776 7524 12782
rect 7472 12718 7524 12724
rect 7484 12442 7512 12718
rect 7472 12436 7524 12442
rect 7472 12378 7524 12384
rect 7380 12300 7432 12306
rect 7380 12242 7432 12248
rect 6920 11756 6972 11762
rect 6920 11698 6972 11704
rect 7576 11694 7604 13126
rect 7716 13084 8024 13093
rect 7716 13082 7722 13084
rect 7778 13082 7802 13084
rect 7858 13082 7882 13084
rect 7938 13082 7962 13084
rect 8018 13082 8024 13084
rect 7778 13030 7780 13082
rect 7960 13030 7962 13082
rect 7716 13028 7722 13030
rect 7778 13028 7802 13030
rect 7858 13028 7882 13030
rect 7938 13028 7962 13030
rect 8018 13028 8024 13030
rect 7716 13019 8024 13028
rect 8128 12306 8156 13330
rect 8116 12300 8168 12306
rect 8116 12242 8168 12248
rect 8220 12238 8248 15150
rect 8300 15156 8352 15162
rect 8300 15098 8352 15104
rect 8312 14414 8340 15098
rect 8404 15094 8432 16526
rect 8496 15502 8524 17478
rect 8484 15496 8536 15502
rect 8484 15438 8536 15444
rect 8392 15088 8444 15094
rect 8392 15030 8444 15036
rect 8300 14408 8352 14414
rect 8300 14350 8352 14356
rect 8404 14074 8432 15030
rect 8496 14414 8524 15438
rect 8484 14408 8536 14414
rect 8484 14350 8536 14356
rect 8392 14068 8444 14074
rect 8392 14010 8444 14016
rect 8404 12866 8432 14010
rect 8588 13394 8616 17478
rect 8680 14550 8708 17478
rect 8956 17462 9076 17490
rect 8944 17332 8996 17338
rect 8944 17274 8996 17280
rect 8956 16590 8984 17274
rect 9048 16590 9076 17462
rect 9140 17338 9168 17614
rect 9416 17542 9444 17682
rect 9220 17536 9272 17542
rect 9220 17478 9272 17484
rect 9404 17536 9456 17542
rect 9404 17478 9456 17484
rect 9496 17536 9548 17542
rect 9496 17478 9548 17484
rect 9128 17332 9180 17338
rect 9128 17274 9180 17280
rect 9232 17134 9260 17478
rect 9312 17332 9364 17338
rect 9312 17274 9364 17280
rect 9220 17128 9272 17134
rect 9220 17070 9272 17076
rect 9128 16992 9180 16998
rect 9128 16934 9180 16940
rect 8944 16584 8996 16590
rect 8944 16526 8996 16532
rect 9036 16584 9088 16590
rect 9036 16526 9088 16532
rect 9140 15484 9168 16934
rect 9232 16794 9260 17070
rect 9220 16788 9272 16794
rect 9220 16730 9272 16736
rect 9324 16590 9352 17274
rect 9416 17202 9444 17478
rect 9404 17196 9456 17202
rect 9404 17138 9456 17144
rect 9508 16658 9536 17478
rect 9600 17202 9628 17818
rect 9692 17762 9720 19860
rect 9692 17734 9812 17762
rect 9784 17678 9812 17734
rect 10980 17678 11008 19860
rect 11127 17980 11435 17989
rect 11127 17978 11133 17980
rect 11189 17978 11213 17980
rect 11269 17978 11293 17980
rect 11349 17978 11373 17980
rect 11429 17978 11435 17980
rect 11189 17926 11191 17978
rect 11371 17926 11373 17978
rect 11127 17924 11133 17926
rect 11189 17924 11213 17926
rect 11269 17924 11293 17926
rect 11349 17924 11373 17926
rect 11429 17924 11435 17926
rect 11127 17915 11435 17924
rect 12268 17678 12296 19860
rect 15198 17980 15506 17989
rect 15198 17978 15204 17980
rect 15260 17978 15284 17980
rect 15340 17978 15364 17980
rect 15420 17978 15444 17980
rect 15500 17978 15506 17980
rect 15260 17926 15262 17978
rect 15442 17926 15444 17978
rect 15198 17924 15204 17926
rect 15260 17924 15284 17926
rect 15340 17924 15364 17926
rect 15420 17924 15444 17926
rect 15500 17924 15506 17926
rect 15198 17915 15506 17924
rect 12348 17876 12400 17882
rect 12348 17818 12400 17824
rect 9772 17672 9824 17678
rect 9772 17614 9824 17620
rect 10968 17672 11020 17678
rect 10968 17614 11020 17620
rect 12256 17672 12308 17678
rect 12256 17614 12308 17620
rect 10048 17604 10100 17610
rect 10048 17546 10100 17552
rect 9588 17196 9640 17202
rect 9588 17138 9640 17144
rect 9600 16998 9628 17138
rect 9864 17128 9916 17134
rect 9864 17070 9916 17076
rect 9588 16992 9640 16998
rect 9588 16934 9640 16940
rect 9876 16794 9904 17070
rect 9864 16788 9916 16794
rect 9864 16730 9916 16736
rect 10060 16726 10088 17546
rect 11520 17536 11572 17542
rect 11520 17478 11572 17484
rect 10876 17128 10928 17134
rect 10876 17070 10928 17076
rect 10324 16992 10376 16998
rect 10324 16934 10376 16940
rect 10048 16720 10100 16726
rect 10048 16662 10100 16668
rect 9496 16652 9548 16658
rect 9496 16594 9548 16600
rect 9312 16584 9364 16590
rect 9312 16526 9364 16532
rect 9312 15496 9364 15502
rect 9140 15456 9312 15484
rect 9312 15438 9364 15444
rect 8668 14544 8720 14550
rect 8668 14486 8720 14492
rect 8680 14278 8708 14486
rect 8668 14272 8720 14278
rect 8668 14214 8720 14220
rect 8576 13388 8628 13394
rect 8576 13330 8628 13336
rect 8588 13002 8616 13330
rect 8944 13252 8996 13258
rect 8944 13194 8996 13200
rect 8588 12974 8708 13002
rect 8956 12986 8984 13194
rect 8484 12912 8536 12918
rect 8404 12860 8484 12866
rect 8404 12854 8536 12860
rect 8404 12838 8524 12854
rect 8208 12232 8260 12238
rect 8208 12174 8260 12180
rect 7716 11996 8024 12005
rect 7716 11994 7722 11996
rect 7778 11994 7802 11996
rect 7858 11994 7882 11996
rect 7938 11994 7962 11996
rect 8018 11994 8024 11996
rect 7778 11942 7780 11994
rect 7960 11942 7962 11994
rect 7716 11940 7722 11942
rect 7778 11940 7802 11942
rect 7858 11940 7882 11942
rect 7938 11940 7962 11942
rect 8018 11940 8024 11942
rect 7716 11931 8024 11940
rect 8220 11762 8248 12174
rect 8208 11756 8260 11762
rect 8208 11698 8260 11704
rect 7564 11688 7616 11694
rect 7564 11630 7616 11636
rect 6920 11552 6972 11558
rect 6920 11494 6972 11500
rect 6932 11286 6960 11494
rect 7056 11452 7364 11461
rect 7056 11450 7062 11452
rect 7118 11450 7142 11452
rect 7198 11450 7222 11452
rect 7278 11450 7302 11452
rect 7358 11450 7364 11452
rect 7118 11398 7120 11450
rect 7300 11398 7302 11450
rect 7056 11396 7062 11398
rect 7118 11396 7142 11398
rect 7198 11396 7222 11398
rect 7278 11396 7302 11398
rect 7358 11396 7364 11398
rect 7056 11387 7364 11396
rect 6920 11280 6972 11286
rect 6920 11222 6972 11228
rect 8404 11218 8432 12838
rect 8680 12238 8708 12974
rect 8944 12980 8996 12986
rect 8944 12922 8996 12928
rect 8956 12306 8984 12922
rect 9324 12782 9352 15438
rect 9588 15428 9640 15434
rect 9588 15370 9640 15376
rect 9404 15360 9456 15366
rect 9404 15302 9456 15308
rect 9416 15026 9444 15302
rect 9600 15162 9628 15370
rect 9588 15156 9640 15162
rect 9588 15098 9640 15104
rect 9404 15020 9456 15026
rect 9404 14962 9456 14968
rect 10232 14476 10284 14482
rect 10232 14418 10284 14424
rect 10244 14074 10272 14418
rect 10336 14414 10364 16934
rect 10888 15434 10916 17070
rect 11127 16892 11435 16901
rect 11127 16890 11133 16892
rect 11189 16890 11213 16892
rect 11269 16890 11293 16892
rect 11349 16890 11373 16892
rect 11429 16890 11435 16892
rect 11189 16838 11191 16890
rect 11371 16838 11373 16890
rect 11127 16836 11133 16838
rect 11189 16836 11213 16838
rect 11269 16836 11293 16838
rect 11349 16836 11373 16838
rect 11429 16836 11435 16838
rect 11127 16827 11435 16836
rect 11127 15804 11435 15813
rect 11127 15802 11133 15804
rect 11189 15802 11213 15804
rect 11269 15802 11293 15804
rect 11349 15802 11373 15804
rect 11429 15802 11435 15804
rect 11189 15750 11191 15802
rect 11371 15750 11373 15802
rect 11127 15748 11133 15750
rect 11189 15748 11213 15750
rect 11269 15748 11293 15750
rect 11349 15748 11373 15750
rect 11429 15748 11435 15750
rect 11127 15739 11435 15748
rect 10876 15428 10928 15434
rect 10876 15370 10928 15376
rect 10324 14408 10376 14414
rect 10324 14350 10376 14356
rect 10232 14068 10284 14074
rect 10232 14010 10284 14016
rect 10140 13932 10192 13938
rect 10140 13874 10192 13880
rect 10152 13326 10180 13874
rect 10336 13394 10364 14350
rect 10416 13932 10468 13938
rect 10416 13874 10468 13880
rect 10428 13462 10456 13874
rect 10416 13456 10468 13462
rect 10416 13398 10468 13404
rect 10324 13388 10376 13394
rect 10324 13330 10376 13336
rect 10140 13320 10192 13326
rect 10140 13262 10192 13268
rect 9588 13184 9640 13190
rect 9588 13126 9640 13132
rect 9600 12918 9628 13126
rect 10888 12918 10916 15370
rect 11127 14716 11435 14725
rect 11127 14714 11133 14716
rect 11189 14714 11213 14716
rect 11269 14714 11293 14716
rect 11349 14714 11373 14716
rect 11429 14714 11435 14716
rect 11189 14662 11191 14714
rect 11371 14662 11373 14714
rect 11127 14660 11133 14662
rect 11189 14660 11213 14662
rect 11269 14660 11293 14662
rect 11349 14660 11373 14662
rect 11429 14660 11435 14662
rect 11127 14651 11435 14660
rect 11127 13628 11435 13637
rect 11127 13626 11133 13628
rect 11189 13626 11213 13628
rect 11269 13626 11293 13628
rect 11349 13626 11373 13628
rect 11429 13626 11435 13628
rect 11189 13574 11191 13626
rect 11371 13574 11373 13626
rect 11127 13572 11133 13574
rect 11189 13572 11213 13574
rect 11269 13572 11293 13574
rect 11349 13572 11373 13574
rect 11429 13572 11435 13574
rect 11127 13563 11435 13572
rect 11532 13410 11560 17478
rect 11787 17436 12095 17445
rect 11787 17434 11793 17436
rect 11849 17434 11873 17436
rect 11929 17434 11953 17436
rect 12009 17434 12033 17436
rect 12089 17434 12095 17436
rect 11849 17382 11851 17434
rect 12031 17382 12033 17434
rect 11787 17380 11793 17382
rect 11849 17380 11873 17382
rect 11929 17380 11953 17382
rect 12009 17380 12033 17382
rect 12089 17380 12095 17382
rect 11787 17371 12095 17380
rect 12360 16998 12388 17818
rect 13084 17604 13136 17610
rect 13084 17546 13136 17552
rect 12532 17536 12584 17542
rect 12532 17478 12584 17484
rect 12348 16992 12400 16998
rect 12348 16934 12400 16940
rect 11704 16652 11756 16658
rect 11704 16594 11756 16600
rect 11612 16584 11664 16590
rect 11612 16526 11664 16532
rect 11624 15366 11652 16526
rect 11716 15706 11744 16594
rect 11787 16348 12095 16357
rect 11787 16346 11793 16348
rect 11849 16346 11873 16348
rect 11929 16346 11953 16348
rect 12009 16346 12033 16348
rect 12089 16346 12095 16348
rect 11849 16294 11851 16346
rect 12031 16294 12033 16346
rect 11787 16292 11793 16294
rect 11849 16292 11873 16294
rect 11929 16292 11953 16294
rect 12009 16292 12033 16294
rect 12089 16292 12095 16294
rect 11787 16283 12095 16292
rect 11704 15700 11756 15706
rect 11704 15642 11756 15648
rect 11704 15496 11756 15502
rect 11704 15438 11756 15444
rect 11612 15360 11664 15366
rect 11612 15302 11664 15308
rect 11624 14482 11652 15302
rect 11716 14482 11744 15438
rect 12256 15428 12308 15434
rect 12256 15370 12308 15376
rect 12164 15360 12216 15366
rect 12164 15302 12216 15308
rect 11787 15260 12095 15269
rect 11787 15258 11793 15260
rect 11849 15258 11873 15260
rect 11929 15258 11953 15260
rect 12009 15258 12033 15260
rect 12089 15258 12095 15260
rect 11849 15206 11851 15258
rect 12031 15206 12033 15258
rect 11787 15204 11793 15206
rect 11849 15204 11873 15206
rect 11929 15204 11953 15206
rect 12009 15204 12033 15206
rect 12089 15204 12095 15206
rect 11787 15195 12095 15204
rect 11888 14952 11940 14958
rect 11888 14894 11940 14900
rect 11796 14816 11848 14822
rect 11796 14758 11848 14764
rect 11808 14550 11836 14758
rect 11900 14618 11928 14894
rect 11888 14612 11940 14618
rect 11888 14554 11940 14560
rect 11796 14544 11848 14550
rect 11796 14486 11848 14492
rect 11612 14476 11664 14482
rect 11612 14418 11664 14424
rect 11704 14476 11756 14482
rect 11704 14418 11756 14424
rect 11808 14362 11836 14486
rect 12176 14414 12204 15302
rect 12268 14822 12296 15370
rect 12256 14816 12308 14822
rect 12256 14758 12308 14764
rect 12268 14414 12296 14758
rect 12360 14550 12388 16934
rect 12544 15502 12572 17478
rect 12992 17128 13044 17134
rect 12992 17070 13044 17076
rect 13004 16794 13032 17070
rect 12992 16788 13044 16794
rect 12992 16730 13044 16736
rect 12624 15632 12676 15638
rect 12624 15574 12676 15580
rect 12532 15496 12584 15502
rect 12532 15438 12584 15444
rect 12348 14544 12400 14550
rect 12348 14486 12400 14492
rect 12544 14414 12572 15438
rect 11716 14334 11836 14362
rect 12164 14408 12216 14414
rect 12164 14350 12216 14356
rect 12256 14408 12308 14414
rect 12256 14350 12308 14356
rect 12532 14408 12584 14414
rect 12532 14350 12584 14356
rect 12440 14340 12492 14346
rect 11440 13382 11560 13410
rect 11612 13456 11664 13462
rect 11612 13398 11664 13404
rect 11440 13326 11468 13382
rect 11624 13326 11652 13398
rect 11060 13320 11112 13326
rect 11060 13262 11112 13268
rect 11428 13320 11480 13326
rect 11428 13262 11480 13268
rect 11612 13320 11664 13326
rect 11612 13262 11664 13268
rect 10968 13252 11020 13258
rect 10968 13194 11020 13200
rect 10980 12986 11008 13194
rect 10968 12980 11020 12986
rect 10968 12922 11020 12928
rect 9588 12912 9640 12918
rect 9588 12854 9640 12860
rect 10876 12912 10928 12918
rect 10876 12854 10928 12860
rect 9312 12776 9364 12782
rect 9312 12718 9364 12724
rect 8944 12300 8996 12306
rect 8944 12242 8996 12248
rect 8668 12232 8720 12238
rect 8668 12174 8720 12180
rect 8668 12096 8720 12102
rect 8668 12038 8720 12044
rect 8680 11898 8708 12038
rect 8668 11892 8720 11898
rect 8668 11834 8720 11840
rect 9324 11218 9352 12718
rect 10888 12442 10916 12854
rect 11072 12594 11100 13262
rect 11520 12776 11572 12782
rect 11716 12764 11744 14334
rect 12440 14282 12492 14288
rect 11787 14172 12095 14181
rect 11787 14170 11793 14172
rect 11849 14170 11873 14172
rect 11929 14170 11953 14172
rect 12009 14170 12033 14172
rect 12089 14170 12095 14172
rect 11849 14118 11851 14170
rect 12031 14118 12033 14170
rect 11787 14116 11793 14118
rect 11849 14116 11873 14118
rect 11929 14116 11953 14118
rect 12009 14116 12033 14118
rect 12089 14116 12095 14118
rect 11787 14107 12095 14116
rect 12452 13394 12480 14282
rect 12636 13462 12664 15574
rect 13096 15502 13124 17546
rect 15858 17436 16166 17445
rect 15858 17434 15864 17436
rect 15920 17434 15944 17436
rect 16000 17434 16024 17436
rect 16080 17434 16104 17436
rect 16160 17434 16166 17436
rect 15920 17382 15922 17434
rect 16102 17382 16104 17434
rect 15858 17380 15864 17382
rect 15920 17380 15944 17382
rect 16000 17380 16024 17382
rect 16080 17380 16104 17382
rect 16160 17380 16166 17382
rect 15858 17371 16166 17380
rect 15198 16892 15506 16901
rect 15198 16890 15204 16892
rect 15260 16890 15284 16892
rect 15340 16890 15364 16892
rect 15420 16890 15444 16892
rect 15500 16890 15506 16892
rect 15260 16838 15262 16890
rect 15442 16838 15444 16890
rect 15198 16836 15204 16838
rect 15260 16836 15284 16838
rect 15340 16836 15364 16838
rect 15420 16836 15444 16838
rect 15500 16836 15506 16838
rect 15198 16827 15506 16836
rect 15858 16348 16166 16357
rect 15858 16346 15864 16348
rect 15920 16346 15944 16348
rect 16000 16346 16024 16348
rect 16080 16346 16104 16348
rect 16160 16346 16166 16348
rect 15920 16294 15922 16346
rect 16102 16294 16104 16346
rect 15858 16292 15864 16294
rect 15920 16292 15944 16294
rect 16000 16292 16024 16294
rect 16080 16292 16104 16294
rect 16160 16292 16166 16294
rect 15858 16283 16166 16292
rect 15198 15804 15506 15813
rect 15198 15802 15204 15804
rect 15260 15802 15284 15804
rect 15340 15802 15364 15804
rect 15420 15802 15444 15804
rect 15500 15802 15506 15804
rect 15260 15750 15262 15802
rect 15442 15750 15444 15802
rect 15198 15748 15204 15750
rect 15260 15748 15284 15750
rect 15340 15748 15364 15750
rect 15420 15748 15444 15750
rect 15500 15748 15506 15750
rect 15198 15739 15506 15748
rect 14924 15564 14976 15570
rect 14924 15506 14976 15512
rect 13084 15496 13136 15502
rect 13084 15438 13136 15444
rect 14936 15434 14964 15506
rect 16580 15496 16632 15502
rect 16580 15438 16632 15444
rect 17040 15496 17092 15502
rect 17040 15438 17092 15444
rect 14924 15428 14976 15434
rect 14924 15370 14976 15376
rect 13268 15360 13320 15366
rect 13268 15302 13320 15308
rect 14188 15360 14240 15366
rect 14188 15302 14240 15308
rect 14556 15360 14608 15366
rect 14556 15302 14608 15308
rect 14740 15360 14792 15366
rect 14740 15302 14792 15308
rect 13280 15026 13308 15302
rect 12900 15020 12952 15026
rect 12900 14962 12952 14968
rect 13268 15020 13320 15026
rect 13268 14962 13320 14968
rect 12624 13456 12676 13462
rect 12624 13398 12676 13404
rect 12440 13388 12492 13394
rect 12440 13330 12492 13336
rect 11787 13084 12095 13093
rect 11787 13082 11793 13084
rect 11849 13082 11873 13084
rect 11929 13082 11953 13084
rect 12009 13082 12033 13084
rect 12089 13082 12095 13084
rect 11849 13030 11851 13082
rect 12031 13030 12033 13082
rect 11787 13028 11793 13030
rect 11849 13028 11873 13030
rect 11929 13028 11953 13030
rect 12009 13028 12033 13030
rect 12089 13028 12095 13030
rect 11787 13019 12095 13028
rect 12912 12850 12940 14962
rect 13280 14414 13308 14962
rect 14096 14952 14148 14958
rect 14096 14894 14148 14900
rect 14108 14618 14136 14894
rect 14096 14612 14148 14618
rect 14096 14554 14148 14560
rect 13268 14408 13320 14414
rect 13268 14350 13320 14356
rect 14200 14346 14228 15302
rect 14372 14952 14424 14958
rect 14372 14894 14424 14900
rect 14384 14414 14412 14894
rect 14568 14482 14596 15302
rect 14752 14482 14780 15302
rect 14936 15162 14964 15370
rect 15858 15260 16166 15269
rect 15858 15258 15864 15260
rect 15920 15258 15944 15260
rect 16000 15258 16024 15260
rect 16080 15258 16104 15260
rect 16160 15258 16166 15260
rect 15920 15206 15922 15258
rect 16102 15206 16104 15258
rect 15858 15204 15864 15206
rect 15920 15204 15944 15206
rect 16000 15204 16024 15206
rect 16080 15204 16104 15206
rect 16160 15204 16166 15206
rect 15858 15195 16166 15204
rect 14924 15156 14976 15162
rect 14924 15098 14976 15104
rect 15660 15088 15712 15094
rect 15660 15030 15712 15036
rect 14924 14952 14976 14958
rect 14924 14894 14976 14900
rect 14936 14618 14964 14894
rect 15568 14816 15620 14822
rect 15568 14758 15620 14764
rect 15198 14716 15506 14725
rect 15198 14714 15204 14716
rect 15260 14714 15284 14716
rect 15340 14714 15364 14716
rect 15420 14714 15444 14716
rect 15500 14714 15506 14716
rect 15260 14662 15262 14714
rect 15442 14662 15444 14714
rect 15198 14660 15204 14662
rect 15260 14660 15284 14662
rect 15340 14660 15364 14662
rect 15420 14660 15444 14662
rect 15500 14660 15506 14662
rect 15198 14651 15506 14660
rect 14924 14612 14976 14618
rect 14924 14554 14976 14560
rect 15580 14482 15608 14758
rect 14556 14476 14608 14482
rect 14556 14418 14608 14424
rect 14740 14476 14792 14482
rect 14740 14418 14792 14424
rect 15568 14476 15620 14482
rect 15568 14418 15620 14424
rect 14372 14408 14424 14414
rect 14372 14350 14424 14356
rect 14188 14340 14240 14346
rect 14188 14282 14240 14288
rect 14280 14340 14332 14346
rect 14280 14282 14332 14288
rect 14292 13870 14320 14282
rect 14384 14074 14412 14350
rect 15672 14346 15700 15030
rect 15660 14340 15712 14346
rect 15660 14282 15712 14288
rect 14372 14068 14424 14074
rect 14372 14010 14424 14016
rect 15672 14006 15700 14282
rect 15858 14172 16166 14181
rect 15858 14170 15864 14172
rect 15920 14170 15944 14172
rect 16000 14170 16024 14172
rect 16080 14170 16104 14172
rect 16160 14170 16166 14172
rect 15920 14118 15922 14170
rect 16102 14118 16104 14170
rect 15858 14116 15864 14118
rect 15920 14116 15944 14118
rect 16000 14116 16024 14118
rect 16080 14116 16104 14118
rect 16160 14116 16166 14118
rect 15858 14107 16166 14116
rect 16592 14074 16620 15438
rect 16856 15360 16908 15366
rect 16856 15302 16908 15308
rect 16868 15065 16896 15302
rect 16854 15056 16910 15065
rect 16854 14991 16910 15000
rect 17052 14618 17080 15438
rect 17040 14612 17092 14618
rect 17040 14554 17092 14560
rect 17038 14376 17094 14385
rect 17038 14311 17094 14320
rect 16580 14068 16632 14074
rect 16580 14010 16632 14016
rect 15660 14000 15712 14006
rect 15660 13942 15712 13948
rect 14280 13864 14332 13870
rect 14280 13806 14332 13812
rect 13176 13320 13228 13326
rect 13176 13262 13228 13268
rect 13544 13320 13596 13326
rect 13544 13262 13596 13268
rect 13188 12986 13216 13262
rect 13176 12980 13228 12986
rect 13176 12922 13228 12928
rect 13556 12850 13584 13262
rect 13728 13184 13780 13190
rect 13728 13126 13780 13132
rect 13740 12986 13768 13126
rect 13728 12980 13780 12986
rect 13728 12922 13780 12928
rect 12900 12844 12952 12850
rect 12900 12786 12952 12792
rect 13544 12844 13596 12850
rect 13544 12786 13596 12792
rect 11572 12736 11744 12764
rect 11520 12718 11572 12724
rect 10980 12566 11100 12594
rect 10876 12436 10928 12442
rect 10796 12406 10876 12434
rect 10232 12096 10284 12102
rect 10232 12038 10284 12044
rect 10244 11898 10272 12038
rect 10232 11892 10284 11898
rect 10232 11834 10284 11840
rect 10324 11892 10376 11898
rect 10324 11834 10376 11840
rect 9772 11824 9824 11830
rect 9772 11766 9824 11772
rect 9784 11558 9812 11766
rect 10336 11762 10364 11834
rect 10324 11756 10376 11762
rect 10324 11698 10376 11704
rect 10416 11756 10468 11762
rect 10416 11698 10468 11704
rect 9772 11552 9824 11558
rect 9772 11494 9824 11500
rect 8392 11212 8444 11218
rect 8392 11154 8444 11160
rect 8668 11212 8720 11218
rect 8668 11154 8720 11160
rect 9312 11212 9364 11218
rect 9312 11154 9364 11160
rect 6828 11144 6880 11150
rect 6828 11086 6880 11092
rect 7716 10908 8024 10917
rect 7716 10906 7722 10908
rect 7778 10906 7802 10908
rect 7858 10906 7882 10908
rect 7938 10906 7962 10908
rect 8018 10906 8024 10908
rect 7778 10854 7780 10906
rect 7960 10854 7962 10906
rect 7716 10852 7722 10854
rect 7778 10852 7802 10854
rect 7858 10852 7882 10854
rect 7938 10852 7962 10854
rect 8018 10852 8024 10854
rect 7716 10843 8024 10852
rect 8404 10810 8432 11154
rect 8484 11008 8536 11014
rect 8484 10950 8536 10956
rect 6736 10804 6788 10810
rect 6736 10746 6788 10752
rect 8392 10804 8444 10810
rect 8392 10746 8444 10752
rect 5868 9540 6040 9568
rect 5816 9522 5868 9528
rect 5540 9512 5592 9518
rect 5540 9454 5592 9460
rect 3424 8968 3476 8974
rect 3424 8910 3476 8916
rect 3516 8968 3568 8974
rect 3516 8910 3568 8916
rect 3424 8288 3476 8294
rect 3528 8276 3556 8910
rect 3712 8906 4016 8922
rect 3700 8900 4016 8906
rect 3752 8894 4016 8900
rect 3700 8842 3752 8848
rect 3645 8732 3953 8741
rect 3645 8730 3651 8732
rect 3707 8730 3731 8732
rect 3787 8730 3811 8732
rect 3867 8730 3891 8732
rect 3947 8730 3953 8732
rect 3707 8678 3709 8730
rect 3889 8678 3891 8730
rect 3645 8676 3651 8678
rect 3707 8676 3731 8678
rect 3787 8676 3811 8678
rect 3867 8676 3891 8678
rect 3947 8676 3953 8678
rect 3645 8667 3953 8676
rect 3988 8566 4016 8894
rect 5356 8900 5408 8906
rect 5356 8842 5408 8848
rect 4712 8832 4764 8838
rect 5368 8786 5396 8842
rect 5552 8838 5580 9454
rect 4712 8774 4764 8780
rect 3976 8560 4028 8566
rect 3976 8502 4028 8508
rect 3988 8294 4016 8502
rect 4724 8498 4752 8774
rect 5276 8758 5396 8786
rect 5540 8832 5592 8838
rect 5540 8774 5592 8780
rect 4712 8492 4764 8498
rect 4712 8434 4764 8440
rect 3476 8248 3556 8276
rect 3976 8288 4028 8294
rect 3424 8230 3476 8236
rect 3976 8230 4028 8236
rect 2985 8188 3293 8197
rect 2985 8186 2991 8188
rect 3047 8186 3071 8188
rect 3127 8186 3151 8188
rect 3207 8186 3231 8188
rect 3287 8186 3293 8188
rect 3047 8134 3049 8186
rect 3229 8134 3231 8186
rect 2985 8132 2991 8134
rect 3047 8132 3071 8134
rect 3127 8132 3151 8134
rect 3207 8132 3231 8134
rect 3287 8132 3293 8134
rect 2985 8123 3293 8132
rect 3148 7744 3200 7750
rect 3424 7744 3476 7750
rect 3200 7704 3372 7732
rect 3148 7686 3200 7692
rect 2872 7200 2924 7206
rect 2872 7142 2924 7148
rect 2780 6452 2832 6458
rect 2780 6394 2832 6400
rect 2884 6338 2912 7142
rect 2985 7100 3293 7109
rect 2985 7098 2991 7100
rect 3047 7098 3071 7100
rect 3127 7098 3151 7100
rect 3207 7098 3231 7100
rect 3287 7098 3293 7100
rect 3047 7046 3049 7098
rect 3229 7046 3231 7098
rect 2985 7044 2991 7046
rect 3047 7044 3071 7046
rect 3127 7044 3151 7046
rect 3207 7044 3231 7046
rect 3287 7044 3293 7046
rect 2985 7035 3293 7044
rect 3344 6798 3372 7704
rect 3424 7686 3476 7692
rect 3436 7342 3464 7686
rect 3645 7644 3953 7653
rect 3645 7642 3651 7644
rect 3707 7642 3731 7644
rect 3787 7642 3811 7644
rect 3867 7642 3891 7644
rect 3947 7642 3953 7644
rect 3707 7590 3709 7642
rect 3889 7590 3891 7642
rect 3645 7588 3651 7590
rect 3707 7588 3731 7590
rect 3787 7588 3811 7590
rect 3867 7588 3891 7590
rect 3947 7588 3953 7590
rect 3645 7579 3953 7588
rect 3988 7478 4016 8230
rect 4724 7478 4752 8434
rect 5276 8294 5304 8758
rect 5552 8566 5580 8774
rect 5736 8634 5764 9522
rect 5724 8628 5776 8634
rect 5724 8570 5776 8576
rect 5540 8560 5592 8566
rect 5540 8502 5592 8508
rect 5264 8288 5316 8294
rect 5264 8230 5316 8236
rect 5276 7478 5304 8230
rect 3608 7472 3660 7478
rect 3608 7414 3660 7420
rect 3976 7472 4028 7478
rect 3976 7414 4028 7420
rect 4712 7472 4764 7478
rect 4712 7414 4764 7420
rect 5264 7472 5316 7478
rect 5264 7414 5316 7420
rect 3424 7336 3476 7342
rect 3424 7278 3476 7284
rect 3332 6792 3384 6798
rect 3332 6734 3384 6740
rect 3436 6662 3464 7278
rect 3620 6730 3648 7414
rect 4068 7336 4120 7342
rect 4068 7278 4120 7284
rect 3976 7200 4028 7206
rect 3976 7142 4028 7148
rect 3988 6798 4016 7142
rect 4080 7002 4108 7278
rect 4068 6996 4120 7002
rect 4068 6938 4120 6944
rect 4066 6896 4122 6905
rect 4066 6831 4122 6840
rect 4080 6798 4108 6831
rect 3976 6792 4028 6798
rect 3976 6734 4028 6740
rect 4068 6792 4120 6798
rect 4068 6734 4120 6740
rect 3608 6724 3660 6730
rect 3528 6684 3608 6712
rect 3424 6656 3476 6662
rect 3424 6598 3476 6604
rect 2504 6316 2556 6322
rect 2504 6258 2556 6264
rect 2792 6310 2912 6338
rect 2516 5846 2544 6258
rect 2504 5840 2556 5846
rect 2504 5782 2556 5788
rect 2516 5710 2544 5782
rect 2792 5710 2820 6310
rect 2872 6248 2924 6254
rect 2872 6190 2924 6196
rect 2412 5704 2464 5710
rect 2412 5646 2464 5652
rect 2504 5704 2556 5710
rect 2504 5646 2556 5652
rect 2780 5704 2832 5710
rect 2780 5646 2832 5652
rect 2884 5642 2912 6190
rect 3332 6112 3384 6118
rect 3332 6054 3384 6060
rect 2985 6012 3293 6021
rect 2985 6010 2991 6012
rect 3047 6010 3071 6012
rect 3127 6010 3151 6012
rect 3207 6010 3231 6012
rect 3287 6010 3293 6012
rect 3047 5958 3049 6010
rect 3229 5958 3231 6010
rect 2985 5956 2991 5958
rect 3047 5956 3071 5958
rect 3127 5956 3151 5958
rect 3207 5956 3231 5958
rect 3287 5956 3293 5958
rect 2985 5947 3293 5956
rect 3148 5908 3200 5914
rect 3148 5850 3200 5856
rect 2872 5636 2924 5642
rect 2872 5578 2924 5584
rect 2780 5568 2832 5574
rect 2780 5510 2832 5516
rect 2792 5370 2820 5510
rect 2780 5364 2832 5370
rect 2780 5306 2832 5312
rect 3160 5302 3188 5850
rect 3344 5778 3372 6054
rect 3528 5914 3556 6684
rect 3608 6666 3660 6672
rect 5080 6656 5132 6662
rect 5080 6598 5132 6604
rect 3645 6556 3953 6565
rect 3645 6554 3651 6556
rect 3707 6554 3731 6556
rect 3787 6554 3811 6556
rect 3867 6554 3891 6556
rect 3947 6554 3953 6556
rect 3707 6502 3709 6554
rect 3889 6502 3891 6554
rect 3645 6500 3651 6502
rect 3707 6500 3731 6502
rect 3787 6500 3811 6502
rect 3867 6500 3891 6502
rect 3947 6500 3953 6502
rect 3645 6491 3953 6500
rect 5092 6458 5120 6598
rect 5080 6452 5132 6458
rect 5080 6394 5132 6400
rect 3516 5908 3568 5914
rect 3516 5850 3568 5856
rect 3332 5772 3384 5778
rect 3332 5714 3384 5720
rect 3424 5772 3476 5778
rect 3424 5714 3476 5720
rect 3516 5772 3568 5778
rect 3516 5714 3568 5720
rect 3240 5636 3292 5642
rect 3240 5578 3292 5584
rect 3148 5296 3200 5302
rect 3148 5238 3200 5244
rect 1584 5160 1636 5166
rect 1584 5102 1636 5108
rect 3252 5114 3280 5578
rect 3344 5302 3372 5714
rect 3332 5296 3384 5302
rect 3332 5238 3384 5244
rect 3436 5234 3464 5714
rect 3528 5370 3556 5714
rect 5092 5642 5120 6394
rect 5080 5636 5132 5642
rect 5080 5578 5132 5584
rect 4528 5568 4580 5574
rect 4528 5510 4580 5516
rect 3645 5468 3953 5477
rect 3645 5466 3651 5468
rect 3707 5466 3731 5468
rect 3787 5466 3811 5468
rect 3867 5466 3891 5468
rect 3947 5466 3953 5468
rect 3707 5414 3709 5466
rect 3889 5414 3891 5466
rect 3645 5412 3651 5414
rect 3707 5412 3731 5414
rect 3787 5412 3811 5414
rect 3867 5412 3891 5414
rect 3947 5412 3953 5414
rect 3645 5403 3953 5412
rect 3516 5364 3568 5370
rect 3516 5306 3568 5312
rect 4540 5302 4568 5510
rect 4528 5296 4580 5302
rect 4528 5238 4580 5244
rect 5092 5250 5120 5578
rect 5276 5302 5304 7414
rect 5828 6662 5856 9522
rect 6368 9376 6420 9382
rect 6368 9318 6420 9324
rect 6380 8974 6408 9318
rect 6184 8968 6236 8974
rect 6184 8910 6236 8916
rect 6368 8968 6420 8974
rect 6368 8910 6420 8916
rect 6552 8968 6604 8974
rect 6552 8910 6604 8916
rect 6196 8498 6224 8910
rect 6460 8832 6512 8838
rect 6460 8774 6512 8780
rect 6184 8492 6236 8498
rect 6184 8434 6236 8440
rect 6196 7546 6224 8434
rect 6472 8430 6500 8774
rect 6564 8634 6592 8910
rect 6552 8628 6604 8634
rect 6552 8570 6604 8576
rect 6748 8498 6776 10746
rect 8496 10742 8524 10950
rect 8484 10736 8536 10742
rect 8484 10678 8536 10684
rect 7564 10668 7616 10674
rect 7564 10610 7616 10616
rect 7056 10364 7364 10373
rect 7056 10362 7062 10364
rect 7118 10362 7142 10364
rect 7198 10362 7222 10364
rect 7278 10362 7302 10364
rect 7358 10362 7364 10364
rect 7118 10310 7120 10362
rect 7300 10310 7302 10362
rect 7056 10308 7062 10310
rect 7118 10308 7142 10310
rect 7198 10308 7222 10310
rect 7278 10308 7302 10310
rect 7358 10308 7364 10310
rect 7056 10299 7364 10308
rect 7380 9512 7432 9518
rect 7380 9454 7432 9460
rect 6920 9376 6972 9382
rect 6920 9318 6972 9324
rect 6932 9042 6960 9318
rect 7056 9276 7364 9285
rect 7056 9274 7062 9276
rect 7118 9274 7142 9276
rect 7198 9274 7222 9276
rect 7278 9274 7302 9276
rect 7358 9274 7364 9276
rect 7118 9222 7120 9274
rect 7300 9222 7302 9274
rect 7056 9220 7062 9222
rect 7118 9220 7142 9222
rect 7198 9220 7222 9222
rect 7278 9220 7302 9222
rect 7358 9220 7364 9222
rect 7056 9211 7364 9220
rect 7392 9178 7420 9454
rect 7380 9172 7432 9178
rect 7432 9132 7512 9160
rect 7380 9114 7432 9120
rect 6920 9036 6972 9042
rect 6920 8978 6972 8984
rect 7380 8900 7432 8906
rect 7380 8842 7432 8848
rect 6736 8492 6788 8498
rect 6736 8434 6788 8440
rect 6460 8424 6512 8430
rect 6460 8366 6512 8372
rect 6920 8424 6972 8430
rect 6920 8366 6972 8372
rect 6932 7818 6960 8366
rect 7056 8188 7364 8197
rect 7056 8186 7062 8188
rect 7118 8186 7142 8188
rect 7198 8186 7222 8188
rect 7278 8186 7302 8188
rect 7358 8186 7364 8188
rect 7118 8134 7120 8186
rect 7300 8134 7302 8186
rect 7056 8132 7062 8134
rect 7118 8132 7142 8134
rect 7198 8132 7222 8134
rect 7278 8132 7302 8134
rect 7358 8132 7364 8134
rect 7056 8123 7364 8132
rect 6920 7812 6972 7818
rect 6920 7754 6972 7760
rect 6932 7562 6960 7754
rect 7392 7562 7420 8842
rect 6184 7540 6236 7546
rect 6184 7482 6236 7488
rect 6840 7534 6960 7562
rect 7300 7546 7420 7562
rect 7300 7540 7432 7546
rect 7300 7534 7380 7540
rect 6840 6746 6868 7534
rect 7300 7478 7328 7534
rect 7380 7482 7432 7488
rect 6920 7472 6972 7478
rect 6920 7414 6972 7420
rect 7288 7472 7340 7478
rect 7484 7426 7512 9132
rect 7576 8430 7604 10610
rect 8208 10464 8260 10470
rect 8208 10406 8260 10412
rect 8116 10056 8168 10062
rect 8116 9998 8168 10004
rect 7716 9820 8024 9829
rect 7716 9818 7722 9820
rect 7778 9818 7802 9820
rect 7858 9818 7882 9820
rect 7938 9818 7962 9820
rect 8018 9818 8024 9820
rect 7778 9766 7780 9818
rect 7960 9766 7962 9818
rect 7716 9764 7722 9766
rect 7778 9764 7802 9766
rect 7858 9764 7882 9766
rect 7938 9764 7962 9766
rect 8018 9764 8024 9766
rect 7716 9755 8024 9764
rect 8128 9586 8156 9998
rect 8220 9654 8248 10406
rect 8300 10056 8352 10062
rect 8300 9998 8352 10004
rect 8208 9648 8260 9654
rect 8208 9590 8260 9596
rect 8116 9580 8168 9586
rect 8116 9522 8168 9528
rect 7716 8732 8024 8741
rect 7716 8730 7722 8732
rect 7778 8730 7802 8732
rect 7858 8730 7882 8732
rect 7938 8730 7962 8732
rect 8018 8730 8024 8732
rect 7778 8678 7780 8730
rect 7960 8678 7962 8730
rect 7716 8676 7722 8678
rect 7778 8676 7802 8678
rect 7858 8676 7882 8678
rect 7938 8676 7962 8678
rect 8018 8676 8024 8678
rect 7716 8667 8024 8676
rect 8128 8634 8156 9522
rect 8116 8628 8168 8634
rect 8116 8570 8168 8576
rect 7564 8424 7616 8430
rect 7564 8366 7616 8372
rect 8220 8022 8248 9590
rect 8312 9518 8340 9998
rect 8484 9920 8536 9926
rect 8484 9862 8536 9868
rect 8496 9518 8524 9862
rect 8680 9586 8708 11154
rect 9220 11076 9272 11082
rect 9220 11018 9272 11024
rect 9232 10810 9260 11018
rect 9220 10804 9272 10810
rect 9220 10746 9272 10752
rect 9784 10674 9812 11494
rect 8760 10668 8812 10674
rect 8760 10610 8812 10616
rect 9772 10668 9824 10674
rect 10336 10656 10364 11698
rect 10428 10810 10456 11698
rect 10692 11688 10744 11694
rect 10692 11630 10744 11636
rect 10704 11354 10732 11630
rect 10692 11348 10744 11354
rect 10692 11290 10744 11296
rect 10416 10804 10468 10810
rect 10416 10746 10468 10752
rect 10704 10742 10732 11290
rect 10796 11082 10824 12406
rect 10980 12434 11008 12566
rect 11127 12540 11435 12549
rect 11127 12538 11133 12540
rect 11189 12538 11213 12540
rect 11269 12538 11293 12540
rect 11349 12538 11373 12540
rect 11429 12538 11435 12540
rect 11189 12486 11191 12538
rect 11371 12486 11373 12538
rect 11127 12484 11133 12486
rect 11189 12484 11213 12486
rect 11269 12484 11293 12486
rect 11349 12484 11373 12486
rect 11429 12484 11435 12486
rect 11127 12475 11435 12484
rect 10980 12406 11100 12434
rect 10876 12378 10928 12384
rect 11072 12102 11100 12406
rect 11060 12096 11112 12102
rect 11060 12038 11112 12044
rect 11532 11762 11560 12718
rect 12912 12442 12940 12786
rect 12900 12436 12952 12442
rect 12952 12406 13124 12434
rect 12900 12378 12952 12384
rect 11787 11996 12095 12005
rect 11787 11994 11793 11996
rect 11849 11994 11873 11996
rect 11929 11994 11953 11996
rect 12009 11994 12033 11996
rect 12089 11994 12095 11996
rect 11849 11942 11851 11994
rect 12031 11942 12033 11994
rect 11787 11940 11793 11942
rect 11849 11940 11873 11942
rect 11929 11940 11953 11942
rect 12009 11940 12033 11942
rect 12089 11940 12095 11942
rect 11787 11931 12095 11940
rect 13096 11830 13124 12406
rect 13556 12306 13584 12786
rect 13544 12300 13596 12306
rect 13544 12242 13596 12248
rect 13740 12238 13768 12922
rect 14292 12850 14320 13806
rect 15198 13628 15506 13637
rect 15198 13626 15204 13628
rect 15260 13626 15284 13628
rect 15340 13626 15364 13628
rect 15420 13626 15444 13628
rect 15500 13626 15506 13628
rect 15260 13574 15262 13626
rect 15442 13574 15444 13626
rect 15198 13572 15204 13574
rect 15260 13572 15284 13574
rect 15340 13572 15364 13574
rect 15420 13572 15444 13574
rect 15500 13572 15506 13574
rect 15198 13563 15506 13572
rect 15672 12850 15700 13942
rect 17052 13938 17080 14311
rect 17040 13932 17092 13938
rect 17040 13874 17092 13880
rect 16212 13728 16264 13734
rect 16212 13670 16264 13676
rect 15858 13084 16166 13093
rect 15858 13082 15864 13084
rect 15920 13082 15944 13084
rect 16000 13082 16024 13084
rect 16080 13082 16104 13084
rect 16160 13082 16166 13084
rect 15920 13030 15922 13082
rect 16102 13030 16104 13082
rect 15858 13028 15864 13030
rect 15920 13028 15944 13030
rect 16000 13028 16024 13030
rect 16080 13028 16104 13030
rect 16160 13028 16166 13030
rect 15858 13019 16166 13028
rect 14280 12844 14332 12850
rect 14280 12786 14332 12792
rect 15660 12844 15712 12850
rect 15660 12786 15712 12792
rect 13820 12776 13872 12782
rect 13820 12718 13872 12724
rect 13832 12238 13860 12718
rect 13728 12232 13780 12238
rect 13728 12174 13780 12180
rect 13820 12232 13872 12238
rect 13820 12174 13872 12180
rect 13084 11824 13136 11830
rect 13084 11766 13136 11772
rect 13728 11824 13780 11830
rect 13728 11766 13780 11772
rect 11520 11756 11572 11762
rect 11520 11698 11572 11704
rect 11532 11558 11560 11698
rect 13740 11694 13768 11766
rect 11796 11688 11848 11694
rect 11796 11630 11848 11636
rect 13636 11688 13688 11694
rect 13636 11630 13688 11636
rect 13728 11688 13780 11694
rect 13728 11630 13780 11636
rect 10876 11552 10928 11558
rect 10876 11494 10928 11500
rect 11520 11552 11572 11558
rect 11520 11494 11572 11500
rect 10888 11218 10916 11494
rect 11127 11452 11435 11461
rect 11127 11450 11133 11452
rect 11189 11450 11213 11452
rect 11269 11450 11293 11452
rect 11349 11450 11373 11452
rect 11429 11450 11435 11452
rect 11189 11398 11191 11450
rect 11371 11398 11373 11450
rect 11127 11396 11133 11398
rect 11189 11396 11213 11398
rect 11269 11396 11293 11398
rect 11349 11396 11373 11398
rect 11429 11396 11435 11398
rect 11127 11387 11435 11396
rect 11808 11354 11836 11630
rect 13268 11552 13320 11558
rect 13268 11494 13320 11500
rect 11796 11348 11848 11354
rect 11796 11290 11848 11296
rect 10876 11212 10928 11218
rect 10876 11154 10928 11160
rect 12808 11212 12860 11218
rect 12808 11154 12860 11160
rect 10968 11144 11020 11150
rect 10968 11086 11020 11092
rect 12440 11144 12492 11150
rect 12440 11086 12492 11092
rect 10784 11076 10836 11082
rect 10784 11018 10836 11024
rect 10692 10736 10744 10742
rect 10692 10678 10744 10684
rect 10416 10668 10468 10674
rect 10336 10628 10416 10656
rect 9772 10610 9824 10616
rect 10416 10610 10468 10616
rect 8668 9580 8720 9586
rect 8668 9522 8720 9528
rect 8300 9512 8352 9518
rect 8300 9454 8352 9460
rect 8484 9512 8536 9518
rect 8484 9454 8536 9460
rect 8312 9178 8340 9454
rect 8300 9172 8352 9178
rect 8300 9114 8352 9120
rect 8772 8974 8800 10610
rect 10980 10538 11008 11086
rect 11787 10908 12095 10917
rect 11787 10906 11793 10908
rect 11849 10906 11873 10908
rect 11929 10906 11953 10908
rect 12009 10906 12033 10908
rect 12089 10906 12095 10908
rect 11849 10854 11851 10906
rect 12031 10854 12033 10906
rect 11787 10852 11793 10854
rect 11849 10852 11873 10854
rect 11929 10852 11953 10854
rect 12009 10852 12033 10854
rect 12089 10852 12095 10854
rect 11787 10843 12095 10852
rect 12452 10674 12480 11086
rect 12820 10810 12848 11154
rect 13280 11150 13308 11494
rect 13648 11354 13676 11630
rect 13636 11348 13688 11354
rect 13636 11290 13688 11296
rect 14292 11218 14320 12786
rect 14556 12776 14608 12782
rect 14556 12718 14608 12724
rect 14568 12442 14596 12718
rect 15198 12540 15506 12549
rect 15198 12538 15204 12540
rect 15260 12538 15284 12540
rect 15340 12538 15364 12540
rect 15420 12538 15444 12540
rect 15500 12538 15506 12540
rect 15260 12486 15262 12538
rect 15442 12486 15444 12538
rect 15198 12484 15204 12486
rect 15260 12484 15284 12486
rect 15340 12484 15364 12486
rect 15420 12484 15444 12486
rect 15500 12484 15506 12486
rect 15198 12475 15506 12484
rect 14556 12436 14608 12442
rect 14556 12378 14608 12384
rect 15108 12232 15160 12238
rect 15108 12174 15160 12180
rect 15120 11898 15148 12174
rect 15568 12164 15620 12170
rect 15568 12106 15620 12112
rect 15108 11892 15160 11898
rect 15108 11834 15160 11840
rect 14924 11756 14976 11762
rect 14924 11698 14976 11704
rect 14280 11212 14332 11218
rect 14280 11154 14332 11160
rect 13268 11144 13320 11150
rect 13268 11086 13320 11092
rect 14936 10810 14964 11698
rect 15580 11694 15608 12106
rect 15568 11688 15620 11694
rect 15568 11630 15620 11636
rect 15672 11642 15700 12786
rect 16028 12640 16080 12646
rect 16028 12582 16080 12588
rect 16040 12238 16068 12582
rect 16224 12442 16252 13670
rect 17040 13320 17092 13326
rect 17040 13262 17092 13268
rect 17052 13025 17080 13262
rect 17038 13016 17094 13025
rect 17038 12951 17094 12960
rect 16212 12436 16264 12442
rect 16212 12378 16264 12384
rect 15752 12232 15804 12238
rect 15752 12174 15804 12180
rect 16028 12232 16080 12238
rect 16028 12174 16080 12180
rect 15764 11830 15792 12174
rect 16212 12164 16264 12170
rect 16212 12106 16264 12112
rect 15858 11996 16166 12005
rect 15858 11994 15864 11996
rect 15920 11994 15944 11996
rect 16000 11994 16024 11996
rect 16080 11994 16104 11996
rect 16160 11994 16166 11996
rect 15920 11942 15922 11994
rect 16102 11942 16104 11994
rect 15858 11940 15864 11942
rect 15920 11940 15944 11942
rect 16000 11940 16024 11942
rect 16080 11940 16104 11942
rect 16160 11940 16166 11942
rect 15858 11931 16166 11940
rect 15752 11824 15804 11830
rect 15752 11766 15804 11772
rect 16224 11694 16252 12106
rect 16488 11756 16540 11762
rect 16488 11698 16540 11704
rect 16580 11756 16632 11762
rect 16580 11698 16632 11704
rect 16212 11688 16264 11694
rect 15108 11552 15160 11558
rect 15108 11494 15160 11500
rect 15120 11234 15148 11494
rect 15198 11452 15506 11461
rect 15198 11450 15204 11452
rect 15260 11450 15284 11452
rect 15340 11450 15364 11452
rect 15420 11450 15444 11452
rect 15500 11450 15506 11452
rect 15260 11398 15262 11450
rect 15442 11398 15444 11450
rect 15198 11396 15204 11398
rect 15260 11396 15284 11398
rect 15340 11396 15364 11398
rect 15420 11396 15444 11398
rect 15500 11396 15506 11398
rect 15198 11387 15506 11396
rect 15120 11206 15240 11234
rect 12808 10804 12860 10810
rect 12808 10746 12860 10752
rect 14924 10804 14976 10810
rect 14924 10746 14976 10752
rect 15212 10742 15240 11206
rect 15200 10736 15252 10742
rect 15200 10678 15252 10684
rect 12440 10668 12492 10674
rect 12440 10610 12492 10616
rect 13268 10668 13320 10674
rect 13268 10610 13320 10616
rect 12808 10600 12860 10606
rect 12808 10542 12860 10548
rect 10968 10532 11020 10538
rect 10968 10474 11020 10480
rect 11704 10464 11756 10470
rect 11704 10406 11756 10412
rect 11127 10364 11435 10373
rect 11127 10362 11133 10364
rect 11189 10362 11213 10364
rect 11269 10362 11293 10364
rect 11349 10362 11373 10364
rect 11429 10362 11435 10364
rect 11189 10310 11191 10362
rect 11371 10310 11373 10362
rect 11127 10308 11133 10310
rect 11189 10308 11213 10310
rect 11269 10308 11293 10310
rect 11349 10308 11373 10310
rect 11429 10308 11435 10310
rect 11127 10299 11435 10308
rect 11716 10130 11744 10406
rect 11704 10124 11756 10130
rect 11704 10066 11756 10072
rect 11428 10056 11480 10062
rect 11428 9998 11480 10004
rect 9956 9648 10008 9654
rect 9956 9590 10008 9596
rect 9128 9512 9180 9518
rect 9128 9454 9180 9460
rect 8852 9444 8904 9450
rect 8852 9386 8904 9392
rect 8864 8974 8892 9386
rect 9140 9110 9168 9454
rect 9128 9104 9180 9110
rect 9128 9046 9180 9052
rect 8760 8968 8812 8974
rect 8760 8910 8812 8916
rect 8852 8968 8904 8974
rect 8852 8910 8904 8916
rect 8668 8900 8720 8906
rect 8668 8842 8720 8848
rect 8392 8832 8444 8838
rect 8392 8774 8444 8780
rect 8404 8566 8432 8774
rect 8392 8560 8444 8566
rect 8392 8502 8444 8508
rect 8680 8498 8708 8842
rect 8668 8492 8720 8498
rect 8668 8434 8720 8440
rect 8208 8016 8260 8022
rect 8208 7958 8260 7964
rect 8668 8016 8720 8022
rect 8668 7958 8720 7964
rect 8300 7948 8352 7954
rect 8300 7890 8352 7896
rect 8208 7880 8260 7886
rect 8208 7822 8260 7828
rect 8116 7812 8168 7818
rect 8116 7754 8168 7760
rect 7564 7744 7616 7750
rect 7564 7686 7616 7692
rect 7288 7414 7340 7420
rect 6932 6866 6960 7414
rect 7392 7398 7512 7426
rect 7392 7342 7420 7398
rect 7380 7336 7432 7342
rect 7380 7278 7432 7284
rect 7056 7100 7364 7109
rect 7056 7098 7062 7100
rect 7118 7098 7142 7100
rect 7198 7098 7222 7100
rect 7278 7098 7302 7100
rect 7358 7098 7364 7100
rect 7118 7046 7120 7098
rect 7300 7046 7302 7098
rect 7056 7044 7062 7046
rect 7118 7044 7142 7046
rect 7198 7044 7222 7046
rect 7278 7044 7302 7046
rect 7358 7044 7364 7046
rect 7056 7035 7364 7044
rect 6920 6860 6972 6866
rect 6920 6802 6972 6808
rect 6840 6730 6960 6746
rect 6840 6724 6972 6730
rect 6840 6718 6920 6724
rect 6920 6666 6972 6672
rect 5816 6656 5868 6662
rect 5816 6598 5868 6604
rect 6460 6656 6512 6662
rect 6460 6598 6512 6604
rect 6472 6458 6500 6598
rect 6460 6452 6512 6458
rect 6460 6394 6512 6400
rect 6932 5914 6960 6666
rect 7056 6012 7364 6021
rect 7056 6010 7062 6012
rect 7118 6010 7142 6012
rect 7198 6010 7222 6012
rect 7278 6010 7302 6012
rect 7358 6010 7364 6012
rect 7118 5958 7120 6010
rect 7300 5958 7302 6010
rect 7056 5956 7062 5958
rect 7118 5956 7142 5958
rect 7198 5956 7222 5958
rect 7278 5956 7302 5958
rect 7358 5956 7364 5958
rect 7056 5947 7364 5956
rect 6920 5908 6972 5914
rect 6920 5850 6972 5856
rect 7196 5908 7248 5914
rect 7196 5850 7248 5856
rect 7012 5840 7064 5846
rect 7012 5782 7064 5788
rect 6828 5772 6880 5778
rect 6828 5714 6880 5720
rect 6552 5568 6604 5574
rect 6552 5510 6604 5516
rect 5264 5296 5316 5302
rect 3424 5228 3476 5234
rect 5092 5222 5212 5250
rect 5264 5238 5316 5244
rect 3424 5170 3476 5176
rect 4160 5160 4212 5166
rect 3252 5098 3372 5114
rect 4160 5102 4212 5108
rect 5080 5160 5132 5166
rect 5080 5102 5132 5108
rect 3252 5092 3384 5098
rect 3252 5086 3332 5092
rect 3332 5034 3384 5040
rect 2985 4924 3293 4933
rect 2985 4922 2991 4924
rect 3047 4922 3071 4924
rect 3127 4922 3151 4924
rect 3207 4922 3231 4924
rect 3287 4922 3293 4924
rect 3047 4870 3049 4922
rect 3229 4870 3231 4922
rect 2985 4868 2991 4870
rect 3047 4868 3071 4870
rect 3127 4868 3151 4870
rect 3207 4868 3231 4870
rect 3287 4868 3293 4870
rect 2985 4859 3293 4868
rect 3645 4380 3953 4389
rect 3645 4378 3651 4380
rect 3707 4378 3731 4380
rect 3787 4378 3811 4380
rect 3867 4378 3891 4380
rect 3947 4378 3953 4380
rect 3707 4326 3709 4378
rect 3889 4326 3891 4378
rect 3645 4324 3651 4326
rect 3707 4324 3731 4326
rect 3787 4324 3811 4326
rect 3867 4324 3891 4326
rect 3947 4324 3953 4326
rect 3645 4315 3953 4324
rect 2985 3836 3293 3845
rect 2985 3834 2991 3836
rect 3047 3834 3071 3836
rect 3127 3834 3151 3836
rect 3207 3834 3231 3836
rect 3287 3834 3293 3836
rect 3047 3782 3049 3834
rect 3229 3782 3231 3834
rect 2985 3780 2991 3782
rect 3047 3780 3071 3782
rect 3127 3780 3151 3782
rect 3207 3780 3231 3782
rect 3287 3780 3293 3782
rect 2985 3771 3293 3780
rect 4172 3602 4200 5102
rect 5092 4690 5120 5102
rect 5080 4684 5132 4690
rect 5080 4626 5132 4632
rect 5184 4282 5212 5222
rect 5276 4486 5304 5238
rect 6564 5166 6592 5510
rect 6552 5160 6604 5166
rect 6552 5102 6604 5108
rect 6368 5024 6420 5030
rect 6368 4966 6420 4972
rect 6380 4690 6408 4966
rect 6564 4690 6592 5102
rect 6368 4684 6420 4690
rect 6368 4626 6420 4632
rect 6552 4684 6604 4690
rect 6552 4626 6604 4632
rect 5264 4480 5316 4486
rect 5264 4422 5316 4428
rect 5172 4276 5224 4282
rect 5172 4218 5224 4224
rect 5080 4140 5132 4146
rect 5080 4082 5132 4088
rect 4712 3936 4764 3942
rect 4712 3878 4764 3884
rect 4160 3596 4212 3602
rect 4160 3538 4212 3544
rect 4068 3460 4120 3466
rect 4068 3402 4120 3408
rect 3645 3292 3953 3301
rect 3645 3290 3651 3292
rect 3707 3290 3731 3292
rect 3787 3290 3811 3292
rect 3867 3290 3891 3292
rect 3947 3290 3953 3292
rect 3707 3238 3709 3290
rect 3889 3238 3891 3290
rect 3645 3236 3651 3238
rect 3707 3236 3731 3238
rect 3787 3236 3811 3238
rect 3867 3236 3891 3238
rect 3947 3236 3953 3238
rect 3645 3227 3953 3236
rect 4080 3194 4108 3402
rect 4724 3194 4752 3878
rect 5092 3738 5120 4082
rect 5080 3732 5132 3738
rect 5080 3674 5132 3680
rect 5276 3602 5304 4422
rect 5816 4276 5868 4282
rect 5816 4218 5868 4224
rect 5448 4140 5500 4146
rect 5448 4082 5500 4088
rect 5264 3596 5316 3602
rect 5264 3538 5316 3544
rect 5460 3466 5488 4082
rect 5828 3466 5856 4218
rect 5448 3460 5500 3466
rect 5448 3402 5500 3408
rect 5816 3460 5868 3466
rect 5816 3402 5868 3408
rect 6276 3460 6328 3466
rect 6276 3402 6328 3408
rect 4068 3188 4120 3194
rect 4068 3130 4120 3136
rect 4712 3188 4764 3194
rect 4712 3130 4764 3136
rect 4724 3058 4752 3130
rect 4712 3052 4764 3058
rect 4712 2994 4764 3000
rect 5356 2984 5408 2990
rect 5356 2926 5408 2932
rect 5368 2854 5396 2926
rect 5356 2848 5408 2854
rect 5356 2790 5408 2796
rect 2985 2748 3293 2757
rect 2985 2746 2991 2748
rect 3047 2746 3071 2748
rect 3127 2746 3151 2748
rect 3207 2746 3231 2748
rect 3287 2746 3293 2748
rect 3047 2694 3049 2746
rect 3229 2694 3231 2746
rect 2985 2692 2991 2694
rect 3047 2692 3071 2694
rect 3127 2692 3151 2694
rect 3207 2692 3231 2694
rect 3287 2692 3293 2694
rect 2985 2683 3293 2692
rect 5460 2650 5488 3402
rect 6092 3392 6144 3398
rect 6092 3334 6144 3340
rect 5724 3188 5776 3194
rect 5724 3130 5776 3136
rect 5736 3058 5764 3130
rect 6104 3058 6132 3334
rect 6288 3194 6316 3402
rect 6276 3188 6328 3194
rect 6276 3130 6328 3136
rect 5724 3052 5776 3058
rect 5724 2994 5776 3000
rect 6092 3052 6144 3058
rect 6092 2994 6144 3000
rect 6840 2650 6868 5714
rect 6920 5704 6972 5710
rect 6920 5646 6972 5652
rect 6932 4826 6960 5646
rect 7024 5370 7052 5782
rect 7208 5710 7236 5850
rect 7196 5704 7248 5710
rect 7392 5658 7420 7278
rect 7576 6866 7604 7686
rect 7716 7644 8024 7653
rect 7716 7642 7722 7644
rect 7778 7642 7802 7644
rect 7858 7642 7882 7644
rect 7938 7642 7962 7644
rect 8018 7642 8024 7644
rect 7778 7590 7780 7642
rect 7960 7590 7962 7642
rect 7716 7588 7722 7590
rect 7778 7588 7802 7590
rect 7858 7588 7882 7590
rect 7938 7588 7962 7590
rect 8018 7588 8024 7590
rect 7716 7579 8024 7588
rect 8128 7546 8156 7754
rect 7656 7540 7708 7546
rect 7656 7482 7708 7488
rect 8116 7540 8168 7546
rect 8116 7482 8168 7488
rect 7564 6860 7616 6866
rect 7564 6802 7616 6808
rect 7668 6644 7696 7482
rect 8024 7404 8076 7410
rect 8024 7346 8076 7352
rect 7196 5646 7248 5652
rect 7300 5630 7420 5658
rect 7576 6616 7696 6644
rect 8036 6644 8064 7346
rect 8128 6798 8156 7482
rect 8220 7002 8248 7822
rect 8208 6996 8260 7002
rect 8208 6938 8260 6944
rect 8312 6798 8340 7890
rect 8484 7744 8536 7750
rect 8484 7686 8536 7692
rect 8496 7342 8524 7686
rect 8680 7410 8708 7958
rect 9140 7818 9168 9046
rect 9772 8288 9824 8294
rect 9772 8230 9824 8236
rect 9784 7954 9812 8230
rect 9772 7948 9824 7954
rect 9772 7890 9824 7896
rect 9968 7818 9996 9590
rect 11440 9466 11468 9998
rect 12440 9988 12492 9994
rect 12440 9930 12492 9936
rect 11787 9820 12095 9829
rect 11787 9818 11793 9820
rect 11849 9818 11873 9820
rect 11929 9818 11953 9820
rect 12009 9818 12033 9820
rect 12089 9818 12095 9820
rect 11849 9766 11851 9818
rect 12031 9766 12033 9818
rect 11787 9764 11793 9766
rect 11849 9764 11873 9766
rect 11929 9764 11953 9766
rect 12009 9764 12033 9766
rect 12089 9764 12095 9766
rect 11787 9755 12095 9764
rect 11440 9438 11560 9466
rect 10692 9376 10744 9382
rect 10692 9318 10744 9324
rect 10600 9036 10652 9042
rect 10600 8978 10652 8984
rect 10612 8634 10640 8978
rect 10704 8974 10732 9318
rect 11127 9276 11435 9285
rect 11127 9274 11133 9276
rect 11189 9274 11213 9276
rect 11269 9274 11293 9276
rect 11349 9274 11373 9276
rect 11429 9274 11435 9276
rect 11189 9222 11191 9274
rect 11371 9222 11373 9274
rect 11127 9220 11133 9222
rect 11189 9220 11213 9222
rect 11269 9220 11293 9222
rect 11349 9220 11373 9222
rect 11429 9220 11435 9222
rect 11127 9211 11435 9220
rect 10692 8968 10744 8974
rect 10692 8910 10744 8916
rect 10704 8634 10732 8910
rect 11060 8832 11112 8838
rect 11060 8774 11112 8780
rect 10600 8628 10652 8634
rect 10600 8570 10652 8576
rect 10692 8628 10744 8634
rect 10692 8570 10744 8576
rect 11072 8566 11100 8774
rect 11060 8560 11112 8566
rect 11060 8502 11112 8508
rect 11532 8430 11560 9438
rect 11787 8732 12095 8741
rect 11787 8730 11793 8732
rect 11849 8730 11873 8732
rect 11929 8730 11953 8732
rect 12009 8730 12033 8732
rect 12089 8730 12095 8732
rect 11849 8678 11851 8730
rect 12031 8678 12033 8730
rect 11787 8676 11793 8678
rect 11849 8676 11873 8678
rect 11929 8676 11953 8678
rect 12009 8676 12033 8678
rect 12089 8676 12095 8678
rect 11787 8667 12095 8676
rect 12452 8566 12480 9930
rect 12716 9920 12768 9926
rect 12716 9862 12768 9868
rect 12440 8560 12492 8566
rect 12440 8502 12492 8508
rect 10416 8424 10468 8430
rect 10416 8366 10468 8372
rect 11520 8424 11572 8430
rect 11520 8366 11572 8372
rect 9128 7812 9180 7818
rect 9128 7754 9180 7760
rect 9956 7812 10008 7818
rect 9956 7754 10008 7760
rect 8668 7404 8720 7410
rect 8668 7346 8720 7352
rect 9140 7342 9168 7754
rect 8484 7336 8536 7342
rect 8484 7278 8536 7284
rect 9128 7336 9180 7342
rect 9128 7278 9180 7284
rect 8116 6792 8168 6798
rect 8116 6734 8168 6740
rect 8300 6792 8352 6798
rect 8300 6734 8352 6740
rect 8116 6656 8168 6662
rect 8036 6616 8116 6644
rect 7012 5364 7064 5370
rect 7012 5306 7064 5312
rect 7300 5098 7328 5630
rect 7380 5364 7432 5370
rect 7576 5352 7604 6616
rect 8116 6598 8168 6604
rect 7716 6556 8024 6565
rect 7716 6554 7722 6556
rect 7778 6554 7802 6556
rect 7858 6554 7882 6556
rect 7938 6554 7962 6556
rect 8018 6554 8024 6556
rect 7778 6502 7780 6554
rect 7960 6502 7962 6554
rect 7716 6500 7722 6502
rect 7778 6500 7802 6502
rect 7858 6500 7882 6502
rect 7938 6500 7962 6502
rect 8018 6500 8024 6502
rect 7716 6491 8024 6500
rect 7716 5468 8024 5477
rect 7716 5466 7722 5468
rect 7778 5466 7802 5468
rect 7858 5466 7882 5468
rect 7938 5466 7962 5468
rect 8018 5466 8024 5468
rect 7778 5414 7780 5466
rect 7960 5414 7962 5466
rect 7716 5412 7722 5414
rect 7778 5412 7802 5414
rect 7858 5412 7882 5414
rect 7938 5412 7962 5414
rect 8018 5412 8024 5414
rect 7716 5403 8024 5412
rect 7748 5364 7800 5370
rect 7576 5324 7748 5352
rect 7380 5306 7432 5312
rect 7288 5092 7340 5098
rect 7288 5034 7340 5040
rect 7056 4924 7364 4933
rect 7056 4922 7062 4924
rect 7118 4922 7142 4924
rect 7198 4922 7222 4924
rect 7278 4922 7302 4924
rect 7358 4922 7364 4924
rect 7118 4870 7120 4922
rect 7300 4870 7302 4922
rect 7056 4868 7062 4870
rect 7118 4868 7142 4870
rect 7198 4868 7222 4870
rect 7278 4868 7302 4870
rect 7358 4868 7364 4870
rect 7056 4859 7364 4868
rect 6920 4820 6972 4826
rect 6920 4762 6972 4768
rect 7392 4690 7420 5306
rect 7564 5160 7616 5166
rect 7564 5102 7616 5108
rect 7576 4826 7604 5102
rect 7564 4820 7616 4826
rect 7564 4762 7616 4768
rect 7380 4684 7432 4690
rect 7380 4626 7432 4632
rect 7668 4570 7696 5324
rect 7748 5306 7800 5312
rect 7576 4542 7696 4570
rect 7576 4214 7604 4542
rect 7716 4380 8024 4389
rect 7716 4378 7722 4380
rect 7778 4378 7802 4380
rect 7858 4378 7882 4380
rect 7938 4378 7962 4380
rect 8018 4378 8024 4380
rect 7778 4326 7780 4378
rect 7960 4326 7962 4378
rect 7716 4324 7722 4326
rect 7778 4324 7802 4326
rect 7858 4324 7882 4326
rect 7938 4324 7962 4326
rect 8018 4324 8024 4326
rect 7716 4315 8024 4324
rect 7564 4208 7616 4214
rect 7564 4150 7616 4156
rect 7056 3836 7364 3845
rect 7056 3834 7062 3836
rect 7118 3834 7142 3836
rect 7198 3834 7222 3836
rect 7278 3834 7302 3836
rect 7358 3834 7364 3836
rect 7118 3782 7120 3834
rect 7300 3782 7302 3834
rect 7056 3780 7062 3782
rect 7118 3780 7142 3782
rect 7198 3780 7222 3782
rect 7278 3780 7302 3782
rect 7358 3780 7364 3782
rect 7056 3771 7364 3780
rect 7576 3466 7604 4150
rect 8128 3738 8156 6598
rect 8208 6316 8260 6322
rect 8208 6258 8260 6264
rect 8220 5914 8248 6258
rect 8208 5908 8260 5914
rect 8208 5850 8260 5856
rect 8220 5710 8248 5850
rect 8208 5704 8260 5710
rect 8208 5646 8260 5652
rect 8208 5160 8260 5166
rect 8208 5102 8260 5108
rect 8220 4146 8248 5102
rect 8208 4140 8260 4146
rect 8208 4082 8260 4088
rect 8116 3732 8168 3738
rect 8116 3674 8168 3680
rect 8220 3602 8248 4082
rect 8208 3596 8260 3602
rect 8208 3538 8260 3544
rect 7564 3460 7616 3466
rect 7564 3402 7616 3408
rect 7576 3126 7604 3402
rect 7716 3292 8024 3301
rect 7716 3290 7722 3292
rect 7778 3290 7802 3292
rect 7858 3290 7882 3292
rect 7938 3290 7962 3292
rect 8018 3290 8024 3292
rect 7778 3238 7780 3290
rect 7960 3238 7962 3290
rect 7716 3236 7722 3238
rect 7778 3236 7802 3238
rect 7858 3236 7882 3238
rect 7938 3236 7962 3238
rect 8018 3236 8024 3238
rect 7716 3227 8024 3236
rect 7564 3120 7616 3126
rect 7564 3062 7616 3068
rect 8220 3058 8248 3538
rect 8208 3052 8260 3058
rect 8208 2994 8260 3000
rect 7056 2748 7364 2757
rect 7056 2746 7062 2748
rect 7118 2746 7142 2748
rect 7198 2746 7222 2748
rect 7278 2746 7302 2748
rect 7358 2746 7364 2748
rect 7118 2694 7120 2746
rect 7300 2694 7302 2746
rect 7056 2692 7062 2694
rect 7118 2692 7142 2694
rect 7198 2692 7222 2694
rect 7278 2692 7302 2694
rect 7358 2692 7364 2694
rect 7056 2683 7364 2692
rect 8312 2650 8340 6734
rect 9140 6322 9168 7278
rect 9968 6390 9996 7754
rect 10428 7546 10456 8366
rect 10784 8356 10836 8362
rect 10784 8298 10836 8304
rect 10796 8090 10824 8298
rect 11127 8188 11435 8197
rect 11127 8186 11133 8188
rect 11189 8186 11213 8188
rect 11269 8186 11293 8188
rect 11349 8186 11373 8188
rect 11429 8186 11435 8188
rect 11189 8134 11191 8186
rect 11371 8134 11373 8186
rect 11127 8132 11133 8134
rect 11189 8132 11213 8134
rect 11269 8132 11293 8134
rect 11349 8132 11373 8134
rect 11429 8132 11435 8134
rect 11127 8123 11435 8132
rect 10784 8084 10836 8090
rect 10784 8026 10836 8032
rect 10876 7812 10928 7818
rect 10876 7754 10928 7760
rect 10692 7744 10744 7750
rect 10692 7686 10744 7692
rect 10416 7540 10468 7546
rect 10416 7482 10468 7488
rect 10704 7478 10732 7686
rect 10692 7472 10744 7478
rect 10692 7414 10744 7420
rect 10888 7410 10916 7754
rect 10324 7404 10376 7410
rect 10324 7346 10376 7352
rect 10876 7404 10928 7410
rect 10876 7346 10928 7352
rect 10048 6656 10100 6662
rect 10048 6598 10100 6604
rect 9956 6384 10008 6390
rect 9956 6326 10008 6332
rect 9128 6316 9180 6322
rect 9128 6258 9180 6264
rect 9864 6248 9916 6254
rect 9864 6190 9916 6196
rect 9876 5914 9904 6190
rect 9968 5914 9996 6326
rect 10060 6118 10088 6598
rect 10048 6112 10100 6118
rect 10048 6054 10100 6060
rect 9864 5908 9916 5914
rect 9864 5850 9916 5856
rect 9956 5908 10008 5914
rect 9956 5850 10008 5856
rect 8944 4072 8996 4078
rect 8944 4014 8996 4020
rect 8956 3738 8984 4014
rect 10060 4010 10088 6054
rect 10140 5704 10192 5710
rect 10140 5646 10192 5652
rect 10152 5370 10180 5646
rect 10140 5364 10192 5370
rect 10140 5306 10192 5312
rect 10232 4548 10284 4554
rect 10232 4490 10284 4496
rect 10244 4214 10272 4490
rect 10232 4208 10284 4214
rect 10232 4150 10284 4156
rect 10048 4004 10100 4010
rect 10048 3946 10100 3952
rect 9864 3936 9916 3942
rect 9864 3878 9916 3884
rect 8944 3732 8996 3738
rect 8944 3674 8996 3680
rect 9876 3534 9904 3878
rect 10060 3534 10088 3946
rect 9036 3528 9088 3534
rect 9036 3470 9088 3476
rect 9864 3528 9916 3534
rect 9864 3470 9916 3476
rect 10048 3528 10100 3534
rect 10048 3470 10100 3476
rect 10140 3528 10192 3534
rect 10140 3470 10192 3476
rect 8668 3392 8720 3398
rect 8668 3334 8720 3340
rect 8680 2990 8708 3334
rect 9048 3194 9076 3470
rect 9036 3188 9088 3194
rect 9036 3130 9088 3136
rect 8668 2984 8720 2990
rect 8668 2926 8720 2932
rect 10152 2650 10180 3470
rect 10336 2774 10364 7346
rect 11532 7342 11560 8366
rect 11787 7644 12095 7653
rect 11787 7642 11793 7644
rect 11849 7642 11873 7644
rect 11929 7642 11953 7644
rect 12009 7642 12033 7644
rect 12089 7642 12095 7644
rect 11849 7590 11851 7642
rect 12031 7590 12033 7642
rect 11787 7588 11793 7590
rect 11849 7588 11873 7590
rect 11929 7588 11953 7590
rect 12009 7588 12033 7590
rect 12089 7588 12095 7590
rect 11787 7579 12095 7588
rect 12452 7478 12480 8502
rect 12728 7750 12756 9862
rect 12820 9722 12848 10542
rect 13280 10266 13308 10610
rect 14924 10600 14976 10606
rect 14924 10542 14976 10548
rect 13728 10464 13780 10470
rect 13728 10406 13780 10412
rect 13268 10260 13320 10266
rect 13268 10202 13320 10208
rect 13084 10124 13136 10130
rect 13084 10066 13136 10072
rect 12808 9716 12860 9722
rect 12808 9658 12860 9664
rect 13096 9654 13124 10066
rect 13740 10062 13768 10406
rect 14936 10266 14964 10542
rect 15198 10364 15506 10373
rect 15198 10362 15204 10364
rect 15260 10362 15284 10364
rect 15340 10362 15364 10364
rect 15420 10362 15444 10364
rect 15500 10362 15506 10364
rect 15260 10310 15262 10362
rect 15442 10310 15444 10362
rect 15198 10308 15204 10310
rect 15260 10308 15284 10310
rect 15340 10308 15364 10310
rect 15420 10308 15444 10310
rect 15500 10308 15506 10310
rect 15198 10299 15506 10308
rect 15580 10266 15608 11630
rect 15672 11614 15792 11642
rect 16500 11665 16528 11698
rect 16212 11630 16264 11636
rect 16486 11656 16542 11665
rect 15764 11558 15792 11614
rect 15660 11552 15712 11558
rect 15660 11494 15712 11500
rect 15752 11552 15804 11558
rect 15752 11494 15804 11500
rect 15672 11218 15700 11494
rect 15660 11212 15712 11218
rect 15660 11154 15712 11160
rect 15764 11082 15792 11494
rect 15752 11076 15804 11082
rect 15752 11018 15804 11024
rect 15858 10908 16166 10917
rect 15858 10906 15864 10908
rect 15920 10906 15944 10908
rect 16000 10906 16024 10908
rect 16080 10906 16104 10908
rect 16160 10906 16166 10908
rect 15920 10854 15922 10906
rect 16102 10854 16104 10906
rect 15858 10852 15864 10854
rect 15920 10852 15944 10854
rect 16000 10852 16024 10854
rect 16080 10852 16104 10854
rect 16160 10852 16166 10854
rect 15858 10843 16166 10852
rect 16224 10810 16252 11630
rect 16486 11591 16542 11600
rect 16488 11212 16540 11218
rect 16488 11154 16540 11160
rect 16212 10804 16264 10810
rect 16212 10746 16264 10752
rect 16500 10742 16528 11154
rect 16592 11014 16620 11698
rect 17040 11144 17092 11150
rect 17040 11086 17092 11092
rect 16580 11008 16632 11014
rect 16580 10950 16632 10956
rect 16856 11008 16908 11014
rect 17052 10985 17080 11086
rect 16856 10950 16908 10956
rect 17038 10976 17094 10985
rect 16592 10810 16620 10950
rect 16580 10804 16632 10810
rect 16580 10746 16632 10752
rect 16488 10736 16540 10742
rect 16488 10678 16540 10684
rect 14924 10260 14976 10266
rect 14924 10202 14976 10208
rect 15568 10260 15620 10266
rect 15568 10202 15620 10208
rect 15384 10124 15436 10130
rect 15384 10066 15436 10072
rect 13728 10056 13780 10062
rect 13728 9998 13780 10004
rect 13084 9648 13136 9654
rect 13084 9590 13136 9596
rect 13740 9586 13768 9998
rect 15396 9722 15424 10066
rect 16500 10062 16528 10678
rect 15752 10056 15804 10062
rect 15752 9998 15804 10004
rect 16488 10056 16540 10062
rect 16488 9998 16540 10004
rect 15384 9716 15436 9722
rect 15384 9658 15436 9664
rect 12808 9580 12860 9586
rect 12808 9522 12860 9528
rect 13728 9580 13780 9586
rect 13728 9522 13780 9528
rect 12716 7744 12768 7750
rect 12716 7686 12768 7692
rect 12440 7472 12492 7478
rect 12440 7414 12492 7420
rect 11520 7336 11572 7342
rect 11520 7278 11572 7284
rect 11127 7100 11435 7109
rect 11127 7098 11133 7100
rect 11189 7098 11213 7100
rect 11269 7098 11293 7100
rect 11349 7098 11373 7100
rect 11429 7098 11435 7100
rect 11189 7046 11191 7098
rect 11371 7046 11373 7098
rect 11127 7044 11133 7046
rect 11189 7044 11213 7046
rect 11269 7044 11293 7046
rect 11349 7044 11373 7046
rect 11429 7044 11435 7046
rect 11127 7035 11435 7044
rect 10968 6724 11020 6730
rect 10968 6666 11020 6672
rect 10980 6390 11008 6666
rect 10968 6384 11020 6390
rect 10968 6326 11020 6332
rect 10784 6180 10836 6186
rect 10784 6122 10836 6128
rect 10600 6112 10652 6118
rect 10600 6054 10652 6060
rect 10612 5710 10640 6054
rect 10692 5840 10744 5846
rect 10692 5782 10744 5788
rect 10600 5704 10652 5710
rect 10600 5646 10652 5652
rect 10600 5568 10652 5574
rect 10600 5510 10652 5516
rect 10612 5166 10640 5510
rect 10600 5160 10652 5166
rect 10600 5102 10652 5108
rect 10704 3534 10732 5782
rect 10796 5710 10824 6122
rect 10980 5846 11008 6326
rect 11127 6012 11435 6021
rect 11127 6010 11133 6012
rect 11189 6010 11213 6012
rect 11269 6010 11293 6012
rect 11349 6010 11373 6012
rect 11429 6010 11435 6012
rect 11189 5958 11191 6010
rect 11371 5958 11373 6010
rect 11127 5956 11133 5958
rect 11189 5956 11213 5958
rect 11269 5956 11293 5958
rect 11349 5956 11373 5958
rect 11429 5956 11435 5958
rect 11127 5947 11435 5956
rect 10968 5840 11020 5846
rect 10968 5782 11020 5788
rect 11532 5778 11560 7278
rect 11787 6556 12095 6565
rect 11787 6554 11793 6556
rect 11849 6554 11873 6556
rect 11929 6554 11953 6556
rect 12009 6554 12033 6556
rect 12089 6554 12095 6556
rect 11849 6502 11851 6554
rect 12031 6502 12033 6554
rect 11787 6500 11793 6502
rect 11849 6500 11873 6502
rect 11929 6500 11953 6502
rect 12009 6500 12033 6502
rect 12089 6500 12095 6502
rect 11787 6491 12095 6500
rect 11704 6180 11756 6186
rect 11704 6122 11756 6128
rect 11520 5772 11572 5778
rect 11520 5714 11572 5720
rect 10784 5704 10836 5710
rect 10784 5646 10836 5652
rect 11532 5234 11560 5714
rect 11520 5228 11572 5234
rect 11520 5170 11572 5176
rect 11127 4924 11435 4933
rect 11127 4922 11133 4924
rect 11189 4922 11213 4924
rect 11269 4922 11293 4924
rect 11349 4922 11373 4924
rect 11429 4922 11435 4924
rect 11189 4870 11191 4922
rect 11371 4870 11373 4922
rect 11127 4868 11133 4870
rect 11189 4868 11213 4870
rect 11269 4868 11293 4870
rect 11349 4868 11373 4870
rect 11429 4868 11435 4870
rect 11127 4859 11435 4868
rect 11127 3836 11435 3845
rect 11127 3834 11133 3836
rect 11189 3834 11213 3836
rect 11269 3834 11293 3836
rect 11349 3834 11373 3836
rect 11429 3834 11435 3836
rect 11189 3782 11191 3834
rect 11371 3782 11373 3834
rect 11127 3780 11133 3782
rect 11189 3780 11213 3782
rect 11269 3780 11293 3782
rect 11349 3780 11373 3782
rect 11429 3780 11435 3782
rect 11127 3771 11435 3780
rect 11532 3602 11560 5170
rect 11520 3596 11572 3602
rect 11520 3538 11572 3544
rect 10692 3528 10744 3534
rect 10692 3470 10744 3476
rect 11152 3460 11204 3466
rect 11152 3402 11204 3408
rect 11164 3194 11192 3402
rect 11152 3188 11204 3194
rect 11152 3130 11204 3136
rect 11532 3058 11560 3538
rect 11612 3460 11664 3466
rect 11612 3402 11664 3408
rect 11624 3126 11652 3402
rect 11612 3120 11664 3126
rect 11612 3062 11664 3068
rect 11520 3052 11572 3058
rect 11520 2994 11572 3000
rect 11520 2916 11572 2922
rect 11520 2858 11572 2864
rect 10244 2746 10364 2774
rect 11127 2748 11435 2757
rect 11127 2746 11133 2748
rect 11189 2746 11213 2748
rect 11269 2746 11293 2748
rect 11349 2746 11373 2748
rect 11429 2746 11435 2748
rect 10244 2650 10272 2746
rect 11189 2694 11191 2746
rect 11371 2694 11373 2746
rect 11127 2692 11133 2694
rect 11189 2692 11213 2694
rect 11269 2692 11293 2694
rect 11349 2692 11373 2694
rect 11429 2692 11435 2694
rect 11127 2683 11435 2692
rect 5448 2644 5500 2650
rect 5448 2586 5500 2592
rect 6828 2644 6880 2650
rect 6828 2586 6880 2592
rect 8300 2644 8352 2650
rect 8300 2586 8352 2592
rect 10140 2644 10192 2650
rect 10140 2586 10192 2592
rect 10232 2644 10284 2650
rect 10232 2586 10284 2592
rect 11532 2582 11560 2858
rect 11716 2774 11744 6122
rect 12452 5914 12480 7414
rect 12728 6662 12756 7686
rect 12820 6730 12848 9522
rect 15198 9276 15506 9285
rect 15198 9274 15204 9276
rect 15260 9274 15284 9276
rect 15340 9274 15364 9276
rect 15420 9274 15444 9276
rect 15500 9274 15506 9276
rect 15260 9222 15262 9274
rect 15442 9222 15444 9274
rect 15198 9220 15204 9222
rect 15260 9220 15284 9222
rect 15340 9220 15364 9222
rect 15420 9220 15444 9222
rect 15500 9220 15506 9222
rect 15198 9211 15506 9220
rect 15764 9178 15792 9998
rect 16212 9920 16264 9926
rect 16212 9862 16264 9868
rect 15858 9820 16166 9829
rect 15858 9818 15864 9820
rect 15920 9818 15944 9820
rect 16000 9818 16024 9820
rect 16080 9818 16104 9820
rect 16160 9818 16166 9820
rect 15920 9766 15922 9818
rect 16102 9766 16104 9818
rect 15858 9764 15864 9766
rect 15920 9764 15944 9766
rect 16000 9764 16024 9766
rect 16080 9764 16104 9766
rect 16160 9764 16166 9766
rect 15858 9755 16166 9764
rect 16224 9722 16252 9862
rect 16592 9738 16620 10746
rect 16868 10674 16896 10950
rect 17038 10911 17094 10920
rect 16856 10668 16908 10674
rect 16856 10610 16908 10616
rect 17040 10668 17092 10674
rect 17040 10610 17092 10616
rect 16868 10062 16896 10610
rect 16948 10600 17000 10606
rect 16948 10542 17000 10548
rect 16856 10056 16908 10062
rect 16856 9998 16908 10004
rect 16212 9716 16264 9722
rect 16212 9658 16264 9664
rect 16500 9710 16620 9738
rect 15936 9580 15988 9586
rect 15936 9522 15988 9528
rect 15948 9178 15976 9522
rect 16120 9512 16172 9518
rect 16120 9454 16172 9460
rect 15752 9172 15804 9178
rect 15752 9114 15804 9120
rect 15936 9172 15988 9178
rect 15936 9114 15988 9120
rect 16132 9042 16160 9454
rect 16120 9036 16172 9042
rect 16120 8978 16172 8984
rect 14096 8968 14148 8974
rect 14096 8910 14148 8916
rect 13912 8900 13964 8906
rect 13912 8842 13964 8848
rect 13924 8634 13952 8842
rect 13912 8628 13964 8634
rect 13912 8570 13964 8576
rect 14108 8498 14136 8910
rect 15016 8832 15068 8838
rect 15016 8774 15068 8780
rect 15028 8566 15056 8774
rect 15858 8732 16166 8741
rect 15858 8730 15864 8732
rect 15920 8730 15944 8732
rect 16000 8730 16024 8732
rect 16080 8730 16104 8732
rect 16160 8730 16166 8732
rect 15920 8678 15922 8730
rect 16102 8678 16104 8730
rect 15858 8676 15864 8678
rect 15920 8676 15944 8678
rect 16000 8676 16024 8678
rect 16080 8676 16104 8678
rect 16160 8676 16166 8678
rect 15858 8667 16166 8676
rect 15016 8560 15068 8566
rect 15016 8502 15068 8508
rect 13636 8492 13688 8498
rect 13636 8434 13688 8440
rect 14096 8492 14148 8498
rect 14096 8434 14148 8440
rect 14556 8492 14608 8498
rect 14556 8434 14608 8440
rect 13452 8424 13504 8430
rect 13452 8366 13504 8372
rect 13464 8090 13492 8366
rect 13452 8084 13504 8090
rect 13452 8026 13504 8032
rect 13544 7880 13596 7886
rect 13544 7822 13596 7828
rect 13452 7472 13504 7478
rect 13452 7414 13504 7420
rect 13464 6798 13492 7414
rect 13556 7342 13584 7822
rect 13648 7410 13676 8434
rect 14004 7812 14056 7818
rect 14004 7754 14056 7760
rect 14016 7546 14044 7754
rect 14280 7744 14332 7750
rect 14280 7686 14332 7692
rect 14004 7540 14056 7546
rect 14004 7482 14056 7488
rect 14292 7478 14320 7686
rect 14280 7472 14332 7478
rect 14280 7414 14332 7420
rect 13636 7404 13688 7410
rect 13636 7346 13688 7352
rect 13820 7404 13872 7410
rect 13820 7346 13872 7352
rect 13544 7336 13596 7342
rect 13832 7290 13860 7346
rect 13544 7278 13596 7284
rect 13556 7002 13584 7278
rect 13740 7262 13860 7290
rect 13544 6996 13596 7002
rect 13544 6938 13596 6944
rect 13740 6798 13768 7262
rect 14292 6798 14320 7414
rect 14568 7410 14596 8434
rect 15198 8188 15506 8197
rect 15198 8186 15204 8188
rect 15260 8186 15284 8188
rect 15340 8186 15364 8188
rect 15420 8186 15444 8188
rect 15500 8186 15506 8188
rect 15260 8134 15262 8186
rect 15442 8134 15444 8186
rect 15198 8132 15204 8134
rect 15260 8132 15284 8134
rect 15340 8132 15364 8134
rect 15420 8132 15444 8134
rect 15500 8132 15506 8134
rect 15198 8123 15506 8132
rect 15858 7644 16166 7653
rect 15858 7642 15864 7644
rect 15920 7642 15944 7644
rect 16000 7642 16024 7644
rect 16080 7642 16104 7644
rect 16160 7642 16166 7644
rect 15920 7590 15922 7642
rect 16102 7590 16104 7642
rect 15858 7588 15864 7590
rect 15920 7588 15944 7590
rect 16000 7588 16024 7590
rect 16080 7588 16104 7590
rect 16160 7588 16166 7590
rect 15858 7579 16166 7588
rect 16224 7426 16252 9658
rect 16304 9580 16356 9586
rect 16304 9522 16356 9528
rect 16316 8974 16344 9522
rect 16304 8968 16356 8974
rect 16304 8910 16356 8916
rect 16316 8634 16344 8910
rect 16396 8900 16448 8906
rect 16396 8842 16448 8848
rect 16304 8628 16356 8634
rect 16304 8570 16356 8576
rect 16408 8566 16436 8842
rect 16396 8560 16448 8566
rect 16396 8502 16448 8508
rect 16408 7478 16436 8502
rect 14556 7404 14608 7410
rect 14556 7346 14608 7352
rect 16132 7398 16252 7426
rect 16396 7472 16448 7478
rect 16396 7414 16448 7420
rect 13452 6792 13504 6798
rect 13452 6734 13504 6740
rect 13728 6792 13780 6798
rect 13728 6734 13780 6740
rect 14280 6792 14332 6798
rect 14280 6734 14332 6740
rect 12808 6724 12860 6730
rect 12808 6666 12860 6672
rect 12716 6656 12768 6662
rect 12716 6598 12768 6604
rect 12440 5908 12492 5914
rect 12440 5850 12492 5856
rect 12452 5794 12480 5850
rect 12452 5766 12572 5794
rect 12544 5642 12572 5766
rect 12440 5636 12492 5642
rect 12440 5578 12492 5584
rect 12532 5636 12584 5642
rect 12532 5578 12584 5584
rect 11787 5468 12095 5477
rect 11787 5466 11793 5468
rect 11849 5466 11873 5468
rect 11929 5466 11953 5468
rect 12009 5466 12033 5468
rect 12089 5466 12095 5468
rect 11849 5414 11851 5466
rect 12031 5414 12033 5466
rect 11787 5412 11793 5414
rect 11849 5412 11873 5414
rect 11929 5412 11953 5414
rect 12009 5412 12033 5414
rect 12089 5412 12095 5414
rect 11787 5403 12095 5412
rect 12452 5370 12480 5578
rect 12440 5364 12492 5370
rect 12440 5306 12492 5312
rect 12544 5302 12572 5578
rect 12532 5296 12584 5302
rect 12532 5238 12584 5244
rect 11787 4380 12095 4389
rect 11787 4378 11793 4380
rect 11849 4378 11873 4380
rect 11929 4378 11953 4380
rect 12009 4378 12033 4380
rect 12089 4378 12095 4380
rect 11849 4326 11851 4378
rect 12031 4326 12033 4378
rect 11787 4324 11793 4326
rect 11849 4324 11873 4326
rect 11929 4324 11953 4326
rect 12009 4324 12033 4326
rect 12089 4324 12095 4326
rect 11787 4315 12095 4324
rect 12728 4146 12756 6598
rect 13740 6322 13768 6734
rect 14464 6452 14516 6458
rect 14464 6394 14516 6400
rect 13728 6316 13780 6322
rect 13728 6258 13780 6264
rect 13912 6316 13964 6322
rect 13912 6258 13964 6264
rect 12900 5636 12952 5642
rect 12900 5578 12952 5584
rect 12624 4140 12676 4146
rect 12624 4082 12676 4088
rect 12716 4140 12768 4146
rect 12716 4082 12768 4088
rect 12256 3936 12308 3942
rect 12256 3878 12308 3884
rect 11787 3292 12095 3301
rect 11787 3290 11793 3292
rect 11849 3290 11873 3292
rect 11929 3290 11953 3292
rect 12009 3290 12033 3292
rect 12089 3290 12095 3292
rect 11849 3238 11851 3290
rect 12031 3238 12033 3290
rect 11787 3236 11793 3238
rect 11849 3236 11873 3238
rect 11929 3236 11953 3238
rect 12009 3236 12033 3238
rect 12089 3236 12095 3238
rect 11787 3227 12095 3236
rect 12268 3058 12296 3878
rect 12636 3738 12664 4082
rect 12912 3738 12940 5578
rect 12992 4208 13044 4214
rect 12992 4150 13044 4156
rect 12624 3732 12676 3738
rect 12624 3674 12676 3680
rect 12900 3732 12952 3738
rect 12900 3674 12952 3680
rect 12912 3398 12940 3674
rect 13004 3466 13032 4150
rect 13452 4140 13504 4146
rect 13452 4082 13504 4088
rect 13464 3534 13492 4082
rect 13740 3738 13768 6258
rect 13924 5914 13952 6258
rect 14004 6112 14056 6118
rect 14004 6054 14056 6060
rect 13912 5908 13964 5914
rect 13912 5850 13964 5856
rect 14016 5370 14044 6054
rect 14476 5710 14504 6394
rect 14568 6338 14596 7346
rect 15568 7336 15620 7342
rect 15568 7278 15620 7284
rect 15198 7100 15506 7109
rect 15198 7098 15204 7100
rect 15260 7098 15284 7100
rect 15340 7098 15364 7100
rect 15420 7098 15444 7100
rect 15500 7098 15506 7100
rect 15260 7046 15262 7098
rect 15442 7046 15444 7098
rect 15198 7044 15204 7046
rect 15260 7044 15284 7046
rect 15340 7044 15364 7046
rect 15420 7044 15444 7046
rect 15500 7044 15506 7046
rect 15198 7035 15506 7044
rect 15580 6866 15608 7278
rect 15568 6860 15620 6866
rect 15568 6802 15620 6808
rect 15660 6792 15712 6798
rect 15660 6734 15712 6740
rect 14568 6310 14688 6338
rect 14556 6248 14608 6254
rect 14556 6190 14608 6196
rect 14568 5846 14596 6190
rect 14556 5840 14608 5846
rect 14556 5782 14608 5788
rect 14464 5704 14516 5710
rect 14464 5646 14516 5652
rect 14096 5568 14148 5574
rect 14096 5510 14148 5516
rect 14004 5364 14056 5370
rect 14004 5306 14056 5312
rect 14016 4622 14044 5306
rect 14108 5234 14136 5510
rect 14660 5302 14688 6310
rect 15198 6012 15506 6021
rect 15198 6010 15204 6012
rect 15260 6010 15284 6012
rect 15340 6010 15364 6012
rect 15420 6010 15444 6012
rect 15500 6010 15506 6012
rect 15260 5958 15262 6010
rect 15442 5958 15444 6010
rect 15198 5956 15204 5958
rect 15260 5956 15284 5958
rect 15340 5956 15364 5958
rect 15420 5956 15444 5958
rect 15500 5956 15506 5958
rect 15198 5947 15506 5956
rect 15672 5710 15700 6734
rect 15752 6724 15804 6730
rect 15752 6666 15804 6672
rect 15764 6322 15792 6666
rect 16132 6662 16160 7398
rect 16304 7200 16356 7206
rect 16304 7142 16356 7148
rect 16212 6860 16264 6866
rect 16212 6802 16264 6808
rect 16120 6656 16172 6662
rect 16120 6598 16172 6604
rect 15858 6556 16166 6565
rect 15858 6554 15864 6556
rect 15920 6554 15944 6556
rect 16000 6554 16024 6556
rect 16080 6554 16104 6556
rect 16160 6554 16166 6556
rect 15920 6502 15922 6554
rect 16102 6502 16104 6554
rect 15858 6500 15864 6502
rect 15920 6500 15944 6502
rect 16000 6500 16024 6502
rect 16080 6500 16104 6502
rect 16160 6500 16166 6502
rect 15858 6491 16166 6500
rect 16224 6322 16252 6802
rect 16316 6798 16344 7142
rect 16304 6792 16356 6798
rect 16304 6734 16356 6740
rect 16304 6656 16356 6662
rect 16304 6598 16356 6604
rect 15752 6316 15804 6322
rect 15752 6258 15804 6264
rect 16212 6316 16264 6322
rect 16212 6258 16264 6264
rect 15752 6112 15804 6118
rect 15752 6054 15804 6060
rect 15764 5778 15792 6054
rect 15752 5772 15804 5778
rect 15752 5714 15804 5720
rect 15660 5704 15712 5710
rect 15660 5646 15712 5652
rect 15672 5386 15700 5646
rect 15858 5468 16166 5477
rect 15858 5466 15864 5468
rect 15920 5466 15944 5468
rect 16000 5466 16024 5468
rect 16080 5466 16104 5468
rect 16160 5466 16166 5468
rect 15920 5414 15922 5466
rect 16102 5414 16104 5466
rect 15858 5412 15864 5414
rect 15920 5412 15944 5414
rect 16000 5412 16024 5414
rect 16080 5412 16104 5414
rect 16160 5412 16166 5414
rect 15858 5403 16166 5412
rect 15580 5370 15700 5386
rect 15568 5364 15700 5370
rect 15620 5358 15700 5364
rect 15568 5306 15620 5312
rect 14464 5296 14516 5302
rect 14464 5238 14516 5244
rect 14648 5296 14700 5302
rect 14648 5238 14700 5244
rect 14096 5228 14148 5234
rect 14096 5170 14148 5176
rect 14108 4758 14136 5170
rect 14280 5024 14332 5030
rect 14280 4966 14332 4972
rect 14096 4752 14148 4758
rect 14096 4694 14148 4700
rect 14292 4622 14320 4966
rect 14476 4758 14504 5238
rect 14556 5160 14608 5166
rect 14556 5102 14608 5108
rect 15752 5160 15804 5166
rect 15752 5102 15804 5108
rect 14568 4826 14596 5102
rect 15198 4924 15506 4933
rect 15198 4922 15204 4924
rect 15260 4922 15284 4924
rect 15340 4922 15364 4924
rect 15420 4922 15444 4924
rect 15500 4922 15506 4924
rect 15260 4870 15262 4922
rect 15442 4870 15444 4922
rect 15198 4868 15204 4870
rect 15260 4868 15284 4870
rect 15340 4868 15364 4870
rect 15420 4868 15444 4870
rect 15500 4868 15506 4870
rect 15198 4859 15506 4868
rect 14556 4820 14608 4826
rect 14556 4762 14608 4768
rect 14464 4752 14516 4758
rect 14464 4694 14516 4700
rect 14004 4616 14056 4622
rect 14004 4558 14056 4564
rect 14280 4616 14332 4622
rect 14280 4558 14332 4564
rect 14096 3936 14148 3942
rect 14096 3878 14148 3884
rect 13728 3732 13780 3738
rect 13728 3674 13780 3680
rect 13452 3528 13504 3534
rect 13452 3470 13504 3476
rect 12992 3460 13044 3466
rect 12992 3402 13044 3408
rect 12900 3392 12952 3398
rect 12900 3334 12952 3340
rect 13360 3392 13412 3398
rect 13360 3334 13412 3340
rect 13372 3194 13400 3334
rect 13360 3188 13412 3194
rect 13360 3130 13412 3136
rect 12256 3052 12308 3058
rect 12256 2994 12308 3000
rect 11888 2984 11940 2990
rect 11888 2926 11940 2932
rect 11624 2746 11744 2774
rect 11624 2650 11652 2746
rect 11612 2644 11664 2650
rect 11612 2586 11664 2592
rect 11520 2576 11572 2582
rect 11520 2518 11572 2524
rect 11900 2446 11928 2926
rect 11980 2848 12032 2854
rect 11980 2790 12032 2796
rect 11992 2514 12020 2790
rect 13464 2650 13492 3470
rect 13636 3392 13688 3398
rect 13636 3334 13688 3340
rect 13648 3126 13676 3334
rect 14108 3126 14136 3878
rect 14476 3602 14504 4694
rect 15764 4554 15792 5102
rect 15752 4548 15804 4554
rect 15752 4490 15804 4496
rect 15292 4480 15344 4486
rect 15292 4422 15344 4428
rect 15304 4146 15332 4422
rect 15764 4162 15792 4490
rect 15858 4380 16166 4389
rect 15858 4378 15864 4380
rect 15920 4378 15944 4380
rect 16000 4378 16024 4380
rect 16080 4378 16104 4380
rect 16160 4378 16166 4380
rect 15920 4326 15922 4378
rect 16102 4326 16104 4378
rect 15858 4324 15864 4326
rect 15920 4324 15944 4326
rect 16000 4324 16024 4326
rect 16080 4324 16104 4326
rect 16160 4324 16166 4326
rect 15858 4315 16166 4324
rect 15292 4140 15344 4146
rect 15292 4082 15344 4088
rect 15476 4140 15528 4146
rect 15476 4082 15528 4088
rect 15568 4140 15620 4146
rect 15764 4134 15884 4162
rect 15568 4082 15620 4088
rect 15304 3924 15332 4082
rect 15120 3896 15332 3924
rect 15488 3924 15516 4082
rect 15580 4026 15608 4082
rect 15580 3998 15792 4026
rect 15660 3936 15712 3942
rect 15488 3896 15608 3924
rect 15120 3618 15148 3896
rect 15198 3836 15506 3845
rect 15198 3834 15204 3836
rect 15260 3834 15284 3836
rect 15340 3834 15364 3836
rect 15420 3834 15444 3836
rect 15500 3834 15506 3836
rect 15260 3782 15262 3834
rect 15442 3782 15444 3834
rect 15198 3780 15204 3782
rect 15260 3780 15284 3782
rect 15340 3780 15364 3782
rect 15420 3780 15444 3782
rect 15500 3780 15506 3782
rect 15198 3771 15506 3780
rect 14464 3596 14516 3602
rect 15120 3590 15240 3618
rect 14464 3538 14516 3544
rect 13636 3120 13688 3126
rect 13636 3062 13688 3068
rect 14096 3120 14148 3126
rect 14096 3062 14148 3068
rect 14476 3058 14504 3538
rect 14648 3460 14700 3466
rect 14648 3402 14700 3408
rect 14660 3194 14688 3402
rect 14648 3188 14700 3194
rect 14648 3130 14700 3136
rect 15212 3058 15240 3590
rect 15384 3392 15436 3398
rect 15384 3334 15436 3340
rect 14464 3052 14516 3058
rect 14464 2994 14516 3000
rect 15200 3052 15252 3058
rect 15200 2994 15252 3000
rect 15396 2922 15424 3334
rect 15580 2922 15608 3896
rect 15660 3878 15712 3884
rect 15672 3058 15700 3878
rect 15764 3398 15792 3998
rect 15856 3466 15884 4134
rect 16316 3534 16344 6598
rect 16408 5234 16436 7414
rect 16396 5228 16448 5234
rect 16396 5170 16448 5176
rect 16500 4010 16528 9710
rect 16856 9580 16908 9586
rect 16856 9522 16908 9528
rect 16868 8974 16896 9522
rect 16960 8974 16988 10542
rect 17052 10305 17080 10610
rect 17038 10296 17094 10305
rect 17038 10231 17094 10240
rect 16856 8968 16908 8974
rect 16856 8910 16908 8916
rect 16948 8968 17000 8974
rect 16948 8910 17000 8916
rect 17038 8936 17094 8945
rect 16868 8634 16896 8910
rect 16856 8628 16908 8634
rect 16856 8570 16908 8576
rect 16672 7200 16724 7206
rect 16672 7142 16724 7148
rect 16684 6798 16712 7142
rect 16960 7018 16988 8910
rect 17038 8871 17094 8880
rect 17052 8498 17080 8871
rect 17040 8492 17092 8498
rect 17040 8434 17092 8440
rect 17040 7880 17092 7886
rect 17040 7822 17092 7828
rect 17052 7585 17080 7822
rect 17038 7576 17094 7585
rect 17038 7511 17094 7520
rect 17040 7404 17092 7410
rect 17040 7346 17092 7352
rect 16868 6990 16988 7018
rect 16868 6798 16896 6990
rect 17052 6905 17080 7346
rect 17038 6896 17094 6905
rect 17038 6831 17094 6840
rect 16672 6792 16724 6798
rect 16672 6734 16724 6740
rect 16856 6792 16908 6798
rect 16856 6734 16908 6740
rect 16764 5568 16816 5574
rect 16764 5510 16816 5516
rect 16776 4690 16804 5510
rect 16764 4684 16816 4690
rect 16764 4626 16816 4632
rect 16580 4140 16632 4146
rect 16580 4082 16632 4088
rect 16488 4004 16540 4010
rect 16488 3946 16540 3952
rect 16592 3738 16620 4082
rect 16580 3732 16632 3738
rect 16580 3674 16632 3680
rect 16304 3528 16356 3534
rect 16304 3470 16356 3476
rect 15844 3460 15896 3466
rect 15844 3402 15896 3408
rect 15752 3392 15804 3398
rect 15752 3334 15804 3340
rect 15764 3126 15792 3334
rect 15858 3292 16166 3301
rect 15858 3290 15864 3292
rect 15920 3290 15944 3292
rect 16000 3290 16024 3292
rect 16080 3290 16104 3292
rect 16160 3290 16166 3292
rect 15920 3238 15922 3290
rect 16102 3238 16104 3290
rect 15858 3236 15864 3238
rect 15920 3236 15944 3238
rect 16000 3236 16024 3238
rect 16080 3236 16104 3238
rect 16160 3236 16166 3238
rect 15858 3227 16166 3236
rect 16592 3194 16620 3674
rect 16868 3670 16896 6734
rect 17040 5704 17092 5710
rect 17040 5646 17092 5652
rect 17052 5545 17080 5646
rect 17038 5536 17094 5545
rect 17038 5471 17094 5480
rect 16856 3664 16908 3670
rect 16856 3606 16908 3612
rect 17040 3528 17092 3534
rect 17038 3496 17040 3505
rect 17092 3496 17094 3505
rect 17038 3431 17094 3440
rect 16580 3188 16632 3194
rect 16580 3130 16632 3136
rect 15752 3120 15804 3126
rect 15752 3062 15804 3068
rect 15660 3052 15712 3058
rect 15660 2994 15712 3000
rect 17040 3052 17092 3058
rect 17040 2994 17092 3000
rect 15384 2916 15436 2922
rect 15384 2858 15436 2864
rect 15568 2916 15620 2922
rect 15568 2858 15620 2864
rect 17052 2825 17080 2994
rect 17038 2816 17094 2825
rect 15198 2748 15506 2757
rect 17038 2751 17094 2760
rect 15198 2746 15204 2748
rect 15260 2746 15284 2748
rect 15340 2746 15364 2748
rect 15420 2746 15444 2748
rect 15500 2746 15506 2748
rect 15260 2694 15262 2746
rect 15442 2694 15444 2746
rect 15198 2692 15204 2694
rect 15260 2692 15284 2694
rect 15340 2692 15364 2694
rect 15420 2692 15444 2694
rect 15500 2692 15506 2694
rect 15198 2683 15506 2692
rect 13452 2644 13504 2650
rect 13452 2586 13504 2592
rect 11980 2508 12032 2514
rect 11980 2450 12032 2456
rect 5172 2440 5224 2446
rect 5172 2382 5224 2388
rect 7104 2440 7156 2446
rect 7104 2382 7156 2388
rect 8392 2440 8444 2446
rect 8392 2382 8444 2388
rect 9680 2440 9732 2446
rect 9680 2382 9732 2388
rect 10324 2440 10376 2446
rect 10324 2382 10376 2388
rect 10968 2440 11020 2446
rect 10968 2382 11020 2388
rect 11888 2440 11940 2446
rect 11888 2382 11940 2388
rect 12900 2440 12952 2446
rect 12900 2382 12952 2388
rect 3645 2204 3953 2213
rect 3645 2202 3651 2204
rect 3707 2202 3731 2204
rect 3787 2202 3811 2204
rect 3867 2202 3891 2204
rect 3947 2202 3953 2204
rect 3707 2150 3709 2202
rect 3889 2150 3891 2202
rect 3645 2148 3651 2150
rect 3707 2148 3731 2150
rect 3787 2148 3811 2150
rect 3867 2148 3891 2150
rect 3947 2148 3953 2150
rect 3645 2139 3953 2148
rect 5184 800 5212 2382
rect 7116 800 7144 2382
rect 7716 2204 8024 2213
rect 7716 2202 7722 2204
rect 7778 2202 7802 2204
rect 7858 2202 7882 2204
rect 7938 2202 7962 2204
rect 8018 2202 8024 2204
rect 7778 2150 7780 2202
rect 7960 2150 7962 2202
rect 7716 2148 7722 2150
rect 7778 2148 7802 2150
rect 7858 2148 7882 2150
rect 7938 2148 7962 2150
rect 8018 2148 8024 2150
rect 7716 2139 8024 2148
rect 8404 800 8432 2382
rect 9692 800 9720 2382
rect 10336 800 10364 2382
rect 10980 800 11008 2382
rect 11787 2204 12095 2213
rect 11787 2202 11793 2204
rect 11849 2202 11873 2204
rect 11929 2202 11953 2204
rect 12009 2202 12033 2204
rect 12089 2202 12095 2204
rect 11849 2150 11851 2202
rect 12031 2150 12033 2202
rect 11787 2148 11793 2150
rect 11849 2148 11873 2150
rect 11929 2148 11953 2150
rect 12009 2148 12033 2150
rect 12089 2148 12095 2150
rect 11787 2139 12095 2148
rect 12912 800 12940 2382
rect 15858 2204 16166 2213
rect 15858 2202 15864 2204
rect 15920 2202 15944 2204
rect 16000 2202 16024 2204
rect 16080 2202 16104 2204
rect 16160 2202 16166 2204
rect 15920 2150 15922 2202
rect 16102 2150 16104 2202
rect 15858 2148 15864 2150
rect 15920 2148 15944 2150
rect 16000 2148 16024 2150
rect 16080 2148 16104 2150
rect 16160 2148 16166 2150
rect 15858 2139 16166 2148
rect 5170 0 5226 800
rect 7102 0 7158 800
rect 8390 0 8446 800
rect 9678 0 9734 800
rect 10322 0 10378 800
rect 10966 0 11022 800
rect 12898 0 12954 800
<< via2 >>
rect 2991 17978 3047 17980
rect 3071 17978 3127 17980
rect 3151 17978 3207 17980
rect 3231 17978 3287 17980
rect 2991 17926 3037 17978
rect 3037 17926 3047 17978
rect 3071 17926 3101 17978
rect 3101 17926 3113 17978
rect 3113 17926 3127 17978
rect 3151 17926 3165 17978
rect 3165 17926 3177 17978
rect 3177 17926 3207 17978
rect 3231 17926 3241 17978
rect 3241 17926 3287 17978
rect 2991 17924 3047 17926
rect 3071 17924 3127 17926
rect 3151 17924 3207 17926
rect 3231 17924 3287 17926
rect 3651 17434 3707 17436
rect 3731 17434 3787 17436
rect 3811 17434 3867 17436
rect 3891 17434 3947 17436
rect 3651 17382 3697 17434
rect 3697 17382 3707 17434
rect 3731 17382 3761 17434
rect 3761 17382 3773 17434
rect 3773 17382 3787 17434
rect 3811 17382 3825 17434
rect 3825 17382 3837 17434
rect 3837 17382 3867 17434
rect 3891 17382 3901 17434
rect 3901 17382 3947 17434
rect 3651 17380 3707 17382
rect 3731 17380 3787 17382
rect 3811 17380 3867 17382
rect 3891 17380 3947 17382
rect 846 17196 902 17232
rect 846 17176 848 17196
rect 848 17176 900 17196
rect 900 17176 902 17196
rect 2991 16890 3047 16892
rect 3071 16890 3127 16892
rect 3151 16890 3207 16892
rect 3231 16890 3287 16892
rect 2991 16838 3037 16890
rect 3037 16838 3047 16890
rect 3071 16838 3101 16890
rect 3101 16838 3113 16890
rect 3113 16838 3127 16890
rect 3151 16838 3165 16890
rect 3165 16838 3177 16890
rect 3177 16838 3207 16890
rect 3231 16838 3241 16890
rect 3241 16838 3287 16890
rect 2991 16836 3047 16838
rect 3071 16836 3127 16838
rect 3151 16836 3207 16838
rect 3231 16836 3287 16838
rect 1030 15680 1086 15736
rect 2991 15802 3047 15804
rect 3071 15802 3127 15804
rect 3151 15802 3207 15804
rect 3231 15802 3287 15804
rect 2991 15750 3037 15802
rect 3037 15750 3047 15802
rect 3071 15750 3101 15802
rect 3101 15750 3113 15802
rect 3113 15750 3127 15802
rect 3151 15750 3165 15802
rect 3165 15750 3177 15802
rect 3177 15750 3207 15802
rect 3231 15750 3241 15802
rect 3241 15750 3287 15802
rect 2991 15748 3047 15750
rect 3071 15748 3127 15750
rect 3151 15748 3207 15750
rect 3231 15748 3287 15750
rect 1398 13640 1454 13696
rect 846 13096 902 13152
rect 846 10784 902 10840
rect 3651 16346 3707 16348
rect 3731 16346 3787 16348
rect 3811 16346 3867 16348
rect 3891 16346 3947 16348
rect 3651 16294 3697 16346
rect 3697 16294 3707 16346
rect 3731 16294 3761 16346
rect 3761 16294 3773 16346
rect 3773 16294 3787 16346
rect 3811 16294 3825 16346
rect 3825 16294 3837 16346
rect 3837 16294 3867 16346
rect 3891 16294 3901 16346
rect 3901 16294 3947 16346
rect 3651 16292 3707 16294
rect 3731 16292 3787 16294
rect 3811 16292 3867 16294
rect 3891 16292 3947 16294
rect 7062 17978 7118 17980
rect 7142 17978 7198 17980
rect 7222 17978 7278 17980
rect 7302 17978 7358 17980
rect 7062 17926 7108 17978
rect 7108 17926 7118 17978
rect 7142 17926 7172 17978
rect 7172 17926 7184 17978
rect 7184 17926 7198 17978
rect 7222 17926 7236 17978
rect 7236 17926 7248 17978
rect 7248 17926 7278 17978
rect 7302 17926 7312 17978
rect 7312 17926 7358 17978
rect 7062 17924 7118 17926
rect 7142 17924 7198 17926
rect 7222 17924 7278 17926
rect 7302 17924 7358 17926
rect 7722 17434 7778 17436
rect 7802 17434 7858 17436
rect 7882 17434 7938 17436
rect 7962 17434 8018 17436
rect 7722 17382 7768 17434
rect 7768 17382 7778 17434
rect 7802 17382 7832 17434
rect 7832 17382 7844 17434
rect 7844 17382 7858 17434
rect 7882 17382 7896 17434
rect 7896 17382 7908 17434
rect 7908 17382 7938 17434
rect 7962 17382 7972 17434
rect 7972 17382 8018 17434
rect 7722 17380 7778 17382
rect 7802 17380 7858 17382
rect 7882 17380 7938 17382
rect 7962 17380 8018 17382
rect 3651 15258 3707 15260
rect 3731 15258 3787 15260
rect 3811 15258 3867 15260
rect 3891 15258 3947 15260
rect 3651 15206 3697 15258
rect 3697 15206 3707 15258
rect 3731 15206 3761 15258
rect 3761 15206 3773 15258
rect 3773 15206 3787 15258
rect 3811 15206 3825 15258
rect 3825 15206 3837 15258
rect 3837 15206 3867 15258
rect 3891 15206 3901 15258
rect 3901 15206 3947 15258
rect 3651 15204 3707 15206
rect 3731 15204 3787 15206
rect 3811 15204 3867 15206
rect 3891 15204 3947 15206
rect 2991 14714 3047 14716
rect 3071 14714 3127 14716
rect 3151 14714 3207 14716
rect 3231 14714 3287 14716
rect 2991 14662 3037 14714
rect 3037 14662 3047 14714
rect 3071 14662 3101 14714
rect 3101 14662 3113 14714
rect 3113 14662 3127 14714
rect 3151 14662 3165 14714
rect 3165 14662 3177 14714
rect 3177 14662 3207 14714
rect 3231 14662 3241 14714
rect 3241 14662 3287 14714
rect 2991 14660 3047 14662
rect 3071 14660 3127 14662
rect 3151 14660 3207 14662
rect 3231 14660 3287 14662
rect 2991 13626 3047 13628
rect 3071 13626 3127 13628
rect 3151 13626 3207 13628
rect 3231 13626 3287 13628
rect 2991 13574 3037 13626
rect 3037 13574 3047 13626
rect 3071 13574 3101 13626
rect 3101 13574 3113 13626
rect 3113 13574 3127 13626
rect 3151 13574 3165 13626
rect 3165 13574 3177 13626
rect 3177 13574 3207 13626
rect 3231 13574 3241 13626
rect 3241 13574 3287 13626
rect 2991 13572 3047 13574
rect 3071 13572 3127 13574
rect 3151 13572 3207 13574
rect 3231 13572 3287 13574
rect 7062 16890 7118 16892
rect 7142 16890 7198 16892
rect 7222 16890 7278 16892
rect 7302 16890 7358 16892
rect 7062 16838 7108 16890
rect 7108 16838 7118 16890
rect 7142 16838 7172 16890
rect 7172 16838 7184 16890
rect 7184 16838 7198 16890
rect 7222 16838 7236 16890
rect 7236 16838 7248 16890
rect 7248 16838 7278 16890
rect 7302 16838 7312 16890
rect 7312 16838 7358 16890
rect 7062 16836 7118 16838
rect 7142 16836 7198 16838
rect 7222 16836 7278 16838
rect 7302 16836 7358 16838
rect 7722 16346 7778 16348
rect 7802 16346 7858 16348
rect 7882 16346 7938 16348
rect 7962 16346 8018 16348
rect 7722 16294 7768 16346
rect 7768 16294 7778 16346
rect 7802 16294 7832 16346
rect 7832 16294 7844 16346
rect 7844 16294 7858 16346
rect 7882 16294 7896 16346
rect 7896 16294 7908 16346
rect 7908 16294 7938 16346
rect 7962 16294 7972 16346
rect 7972 16294 8018 16346
rect 7722 16292 7778 16294
rect 7802 16292 7858 16294
rect 7882 16292 7938 16294
rect 7962 16292 8018 16294
rect 7062 15802 7118 15804
rect 7142 15802 7198 15804
rect 7222 15802 7278 15804
rect 7302 15802 7358 15804
rect 7062 15750 7108 15802
rect 7108 15750 7118 15802
rect 7142 15750 7172 15802
rect 7172 15750 7184 15802
rect 7184 15750 7198 15802
rect 7222 15750 7236 15802
rect 7236 15750 7248 15802
rect 7248 15750 7278 15802
rect 7302 15750 7312 15802
rect 7312 15750 7358 15802
rect 7062 15748 7118 15750
rect 7142 15748 7198 15750
rect 7222 15748 7278 15750
rect 7302 15748 7358 15750
rect 7062 14714 7118 14716
rect 7142 14714 7198 14716
rect 7222 14714 7278 14716
rect 7302 14714 7358 14716
rect 7062 14662 7108 14714
rect 7108 14662 7118 14714
rect 7142 14662 7172 14714
rect 7172 14662 7184 14714
rect 7184 14662 7198 14714
rect 7222 14662 7236 14714
rect 7236 14662 7248 14714
rect 7248 14662 7278 14714
rect 7302 14662 7312 14714
rect 7312 14662 7358 14714
rect 7062 14660 7118 14662
rect 7142 14660 7198 14662
rect 7222 14660 7278 14662
rect 7302 14660 7358 14662
rect 7722 15258 7778 15260
rect 7802 15258 7858 15260
rect 7882 15258 7938 15260
rect 7962 15258 8018 15260
rect 7722 15206 7768 15258
rect 7768 15206 7778 15258
rect 7802 15206 7832 15258
rect 7832 15206 7844 15258
rect 7844 15206 7858 15258
rect 7882 15206 7896 15258
rect 7896 15206 7908 15258
rect 7908 15206 7938 15258
rect 7962 15206 7972 15258
rect 7972 15206 8018 15258
rect 7722 15204 7778 15206
rect 7802 15204 7858 15206
rect 7882 15204 7938 15206
rect 7962 15204 8018 15206
rect 3651 14170 3707 14172
rect 3731 14170 3787 14172
rect 3811 14170 3867 14172
rect 3891 14170 3947 14172
rect 3651 14118 3697 14170
rect 3697 14118 3707 14170
rect 3731 14118 3761 14170
rect 3761 14118 3773 14170
rect 3773 14118 3787 14170
rect 3811 14118 3825 14170
rect 3825 14118 3837 14170
rect 3837 14118 3867 14170
rect 3891 14118 3901 14170
rect 3901 14118 3947 14170
rect 3651 14116 3707 14118
rect 3731 14116 3787 14118
rect 3811 14116 3867 14118
rect 3891 14116 3947 14118
rect 2991 12538 3047 12540
rect 3071 12538 3127 12540
rect 3151 12538 3207 12540
rect 3231 12538 3287 12540
rect 2991 12486 3037 12538
rect 3037 12486 3047 12538
rect 3071 12486 3101 12538
rect 3101 12486 3113 12538
rect 3113 12486 3127 12538
rect 3151 12486 3165 12538
rect 3165 12486 3177 12538
rect 3177 12486 3207 12538
rect 3231 12486 3241 12538
rect 3241 12486 3287 12538
rect 2991 12484 3047 12486
rect 3071 12484 3127 12486
rect 3151 12484 3207 12486
rect 3231 12484 3287 12486
rect 2991 11450 3047 11452
rect 3071 11450 3127 11452
rect 3151 11450 3207 11452
rect 3231 11450 3287 11452
rect 2991 11398 3037 11450
rect 3037 11398 3047 11450
rect 3071 11398 3101 11450
rect 3101 11398 3113 11450
rect 3113 11398 3127 11450
rect 3151 11398 3165 11450
rect 3165 11398 3177 11450
rect 3177 11398 3207 11450
rect 3231 11398 3241 11450
rect 3241 11398 3287 11450
rect 2991 11396 3047 11398
rect 3071 11396 3127 11398
rect 3151 11396 3207 11398
rect 3231 11396 3287 11398
rect 1398 9560 1454 9616
rect 2991 10362 3047 10364
rect 3071 10362 3127 10364
rect 3151 10362 3207 10364
rect 3231 10362 3287 10364
rect 2991 10310 3037 10362
rect 3037 10310 3047 10362
rect 3071 10310 3101 10362
rect 3101 10310 3113 10362
rect 3113 10310 3127 10362
rect 3151 10310 3165 10362
rect 3165 10310 3177 10362
rect 3177 10310 3207 10362
rect 3231 10310 3241 10362
rect 3241 10310 3287 10362
rect 2991 10308 3047 10310
rect 3071 10308 3127 10310
rect 3151 10308 3207 10310
rect 3231 10308 3287 10310
rect 3651 13082 3707 13084
rect 3731 13082 3787 13084
rect 3811 13082 3867 13084
rect 3891 13082 3947 13084
rect 3651 13030 3697 13082
rect 3697 13030 3707 13082
rect 3731 13030 3761 13082
rect 3761 13030 3773 13082
rect 3773 13030 3787 13082
rect 3811 13030 3825 13082
rect 3825 13030 3837 13082
rect 3837 13030 3867 13082
rect 3891 13030 3901 13082
rect 3901 13030 3947 13082
rect 3651 13028 3707 13030
rect 3731 13028 3787 13030
rect 3811 13028 3867 13030
rect 3891 13028 3947 13030
rect 3651 11994 3707 11996
rect 3731 11994 3787 11996
rect 3811 11994 3867 11996
rect 3891 11994 3947 11996
rect 3651 11942 3697 11994
rect 3697 11942 3707 11994
rect 3731 11942 3761 11994
rect 3761 11942 3773 11994
rect 3773 11942 3787 11994
rect 3811 11942 3825 11994
rect 3825 11942 3837 11994
rect 3837 11942 3867 11994
rect 3891 11942 3901 11994
rect 3901 11942 3947 11994
rect 3651 11940 3707 11942
rect 3731 11940 3787 11942
rect 3811 11940 3867 11942
rect 3891 11940 3947 11942
rect 3651 10906 3707 10908
rect 3731 10906 3787 10908
rect 3811 10906 3867 10908
rect 3891 10906 3947 10908
rect 3651 10854 3697 10906
rect 3697 10854 3707 10906
rect 3731 10854 3761 10906
rect 3761 10854 3773 10906
rect 3773 10854 3787 10906
rect 3811 10854 3825 10906
rect 3825 10854 3837 10906
rect 3837 10854 3867 10906
rect 3891 10854 3901 10906
rect 3901 10854 3947 10906
rect 3651 10852 3707 10854
rect 3731 10852 3787 10854
rect 3811 10852 3867 10854
rect 3891 10852 3947 10854
rect 3651 9818 3707 9820
rect 3731 9818 3787 9820
rect 3811 9818 3867 9820
rect 3891 9818 3947 9820
rect 3651 9766 3697 9818
rect 3697 9766 3707 9818
rect 3731 9766 3761 9818
rect 3761 9766 3773 9818
rect 3773 9766 3787 9818
rect 3811 9766 3825 9818
rect 3825 9766 3837 9818
rect 3837 9766 3867 9818
rect 3891 9766 3901 9818
rect 3901 9766 3947 9818
rect 3651 9764 3707 9766
rect 3731 9764 3787 9766
rect 3811 9764 3867 9766
rect 3891 9764 3947 9766
rect 2962 9580 3018 9616
rect 2962 9560 2964 9580
rect 2964 9560 3016 9580
rect 3016 9560 3018 9580
rect 2410 9460 2412 9480
rect 2412 9460 2464 9480
rect 2464 9460 2466 9480
rect 846 8744 902 8800
rect 846 7656 902 7712
rect 2410 9424 2466 9460
rect 7722 14170 7778 14172
rect 7802 14170 7858 14172
rect 7882 14170 7938 14172
rect 7962 14170 8018 14172
rect 7722 14118 7768 14170
rect 7768 14118 7778 14170
rect 7802 14118 7832 14170
rect 7832 14118 7844 14170
rect 7844 14118 7858 14170
rect 7882 14118 7896 14170
rect 7896 14118 7908 14170
rect 7908 14118 7938 14170
rect 7962 14118 7972 14170
rect 7972 14118 8018 14170
rect 7722 14116 7778 14118
rect 7802 14116 7858 14118
rect 7882 14116 7938 14118
rect 7962 14116 8018 14118
rect 7062 13626 7118 13628
rect 7142 13626 7198 13628
rect 7222 13626 7278 13628
rect 7302 13626 7358 13628
rect 7062 13574 7108 13626
rect 7108 13574 7118 13626
rect 7142 13574 7172 13626
rect 7172 13574 7184 13626
rect 7184 13574 7198 13626
rect 7222 13574 7236 13626
rect 7236 13574 7248 13626
rect 7248 13574 7278 13626
rect 7302 13574 7312 13626
rect 7312 13574 7358 13626
rect 7062 13572 7118 13574
rect 7142 13572 7198 13574
rect 7222 13572 7278 13574
rect 7302 13572 7358 13574
rect 3422 9560 3478 9616
rect 1674 8200 1730 8256
rect 1398 5480 1454 5536
rect 3330 9424 3386 9480
rect 2991 9274 3047 9276
rect 3071 9274 3127 9276
rect 3151 9274 3207 9276
rect 3231 9274 3287 9276
rect 2991 9222 3037 9274
rect 3037 9222 3047 9274
rect 3071 9222 3101 9274
rect 3101 9222 3113 9274
rect 3113 9222 3127 9274
rect 3151 9222 3165 9274
rect 3165 9222 3177 9274
rect 3177 9222 3207 9274
rect 3231 9222 3241 9274
rect 3241 9222 3287 9274
rect 2991 9220 3047 9222
rect 3071 9220 3127 9222
rect 3151 9220 3207 9222
rect 3231 9220 3287 9222
rect 7062 12538 7118 12540
rect 7142 12538 7198 12540
rect 7222 12538 7278 12540
rect 7302 12538 7358 12540
rect 7062 12486 7108 12538
rect 7108 12486 7118 12538
rect 7142 12486 7172 12538
rect 7172 12486 7184 12538
rect 7184 12486 7198 12538
rect 7222 12486 7236 12538
rect 7236 12486 7248 12538
rect 7248 12486 7278 12538
rect 7302 12486 7312 12538
rect 7312 12486 7358 12538
rect 7062 12484 7118 12486
rect 7142 12484 7198 12486
rect 7222 12484 7278 12486
rect 7302 12484 7358 12486
rect 7722 13082 7778 13084
rect 7802 13082 7858 13084
rect 7882 13082 7938 13084
rect 7962 13082 8018 13084
rect 7722 13030 7768 13082
rect 7768 13030 7778 13082
rect 7802 13030 7832 13082
rect 7832 13030 7844 13082
rect 7844 13030 7858 13082
rect 7882 13030 7896 13082
rect 7896 13030 7908 13082
rect 7908 13030 7938 13082
rect 7962 13030 7972 13082
rect 7972 13030 8018 13082
rect 7722 13028 7778 13030
rect 7802 13028 7858 13030
rect 7882 13028 7938 13030
rect 7962 13028 8018 13030
rect 11133 17978 11189 17980
rect 11213 17978 11269 17980
rect 11293 17978 11349 17980
rect 11373 17978 11429 17980
rect 11133 17926 11179 17978
rect 11179 17926 11189 17978
rect 11213 17926 11243 17978
rect 11243 17926 11255 17978
rect 11255 17926 11269 17978
rect 11293 17926 11307 17978
rect 11307 17926 11319 17978
rect 11319 17926 11349 17978
rect 11373 17926 11383 17978
rect 11383 17926 11429 17978
rect 11133 17924 11189 17926
rect 11213 17924 11269 17926
rect 11293 17924 11349 17926
rect 11373 17924 11429 17926
rect 15204 17978 15260 17980
rect 15284 17978 15340 17980
rect 15364 17978 15420 17980
rect 15444 17978 15500 17980
rect 15204 17926 15250 17978
rect 15250 17926 15260 17978
rect 15284 17926 15314 17978
rect 15314 17926 15326 17978
rect 15326 17926 15340 17978
rect 15364 17926 15378 17978
rect 15378 17926 15390 17978
rect 15390 17926 15420 17978
rect 15444 17926 15454 17978
rect 15454 17926 15500 17978
rect 15204 17924 15260 17926
rect 15284 17924 15340 17926
rect 15364 17924 15420 17926
rect 15444 17924 15500 17926
rect 7722 11994 7778 11996
rect 7802 11994 7858 11996
rect 7882 11994 7938 11996
rect 7962 11994 8018 11996
rect 7722 11942 7768 11994
rect 7768 11942 7778 11994
rect 7802 11942 7832 11994
rect 7832 11942 7844 11994
rect 7844 11942 7858 11994
rect 7882 11942 7896 11994
rect 7896 11942 7908 11994
rect 7908 11942 7938 11994
rect 7962 11942 7972 11994
rect 7972 11942 8018 11994
rect 7722 11940 7778 11942
rect 7802 11940 7858 11942
rect 7882 11940 7938 11942
rect 7962 11940 8018 11942
rect 7062 11450 7118 11452
rect 7142 11450 7198 11452
rect 7222 11450 7278 11452
rect 7302 11450 7358 11452
rect 7062 11398 7108 11450
rect 7108 11398 7118 11450
rect 7142 11398 7172 11450
rect 7172 11398 7184 11450
rect 7184 11398 7198 11450
rect 7222 11398 7236 11450
rect 7236 11398 7248 11450
rect 7248 11398 7278 11450
rect 7302 11398 7312 11450
rect 7312 11398 7358 11450
rect 7062 11396 7118 11398
rect 7142 11396 7198 11398
rect 7222 11396 7278 11398
rect 7302 11396 7358 11398
rect 11133 16890 11189 16892
rect 11213 16890 11269 16892
rect 11293 16890 11349 16892
rect 11373 16890 11429 16892
rect 11133 16838 11179 16890
rect 11179 16838 11189 16890
rect 11213 16838 11243 16890
rect 11243 16838 11255 16890
rect 11255 16838 11269 16890
rect 11293 16838 11307 16890
rect 11307 16838 11319 16890
rect 11319 16838 11349 16890
rect 11373 16838 11383 16890
rect 11383 16838 11429 16890
rect 11133 16836 11189 16838
rect 11213 16836 11269 16838
rect 11293 16836 11349 16838
rect 11373 16836 11429 16838
rect 11133 15802 11189 15804
rect 11213 15802 11269 15804
rect 11293 15802 11349 15804
rect 11373 15802 11429 15804
rect 11133 15750 11179 15802
rect 11179 15750 11189 15802
rect 11213 15750 11243 15802
rect 11243 15750 11255 15802
rect 11255 15750 11269 15802
rect 11293 15750 11307 15802
rect 11307 15750 11319 15802
rect 11319 15750 11349 15802
rect 11373 15750 11383 15802
rect 11383 15750 11429 15802
rect 11133 15748 11189 15750
rect 11213 15748 11269 15750
rect 11293 15748 11349 15750
rect 11373 15748 11429 15750
rect 11133 14714 11189 14716
rect 11213 14714 11269 14716
rect 11293 14714 11349 14716
rect 11373 14714 11429 14716
rect 11133 14662 11179 14714
rect 11179 14662 11189 14714
rect 11213 14662 11243 14714
rect 11243 14662 11255 14714
rect 11255 14662 11269 14714
rect 11293 14662 11307 14714
rect 11307 14662 11319 14714
rect 11319 14662 11349 14714
rect 11373 14662 11383 14714
rect 11383 14662 11429 14714
rect 11133 14660 11189 14662
rect 11213 14660 11269 14662
rect 11293 14660 11349 14662
rect 11373 14660 11429 14662
rect 11133 13626 11189 13628
rect 11213 13626 11269 13628
rect 11293 13626 11349 13628
rect 11373 13626 11429 13628
rect 11133 13574 11179 13626
rect 11179 13574 11189 13626
rect 11213 13574 11243 13626
rect 11243 13574 11255 13626
rect 11255 13574 11269 13626
rect 11293 13574 11307 13626
rect 11307 13574 11319 13626
rect 11319 13574 11349 13626
rect 11373 13574 11383 13626
rect 11383 13574 11429 13626
rect 11133 13572 11189 13574
rect 11213 13572 11269 13574
rect 11293 13572 11349 13574
rect 11373 13572 11429 13574
rect 11793 17434 11849 17436
rect 11873 17434 11929 17436
rect 11953 17434 12009 17436
rect 12033 17434 12089 17436
rect 11793 17382 11839 17434
rect 11839 17382 11849 17434
rect 11873 17382 11903 17434
rect 11903 17382 11915 17434
rect 11915 17382 11929 17434
rect 11953 17382 11967 17434
rect 11967 17382 11979 17434
rect 11979 17382 12009 17434
rect 12033 17382 12043 17434
rect 12043 17382 12089 17434
rect 11793 17380 11849 17382
rect 11873 17380 11929 17382
rect 11953 17380 12009 17382
rect 12033 17380 12089 17382
rect 11793 16346 11849 16348
rect 11873 16346 11929 16348
rect 11953 16346 12009 16348
rect 12033 16346 12089 16348
rect 11793 16294 11839 16346
rect 11839 16294 11849 16346
rect 11873 16294 11903 16346
rect 11903 16294 11915 16346
rect 11915 16294 11929 16346
rect 11953 16294 11967 16346
rect 11967 16294 11979 16346
rect 11979 16294 12009 16346
rect 12033 16294 12043 16346
rect 12043 16294 12089 16346
rect 11793 16292 11849 16294
rect 11873 16292 11929 16294
rect 11953 16292 12009 16294
rect 12033 16292 12089 16294
rect 11793 15258 11849 15260
rect 11873 15258 11929 15260
rect 11953 15258 12009 15260
rect 12033 15258 12089 15260
rect 11793 15206 11839 15258
rect 11839 15206 11849 15258
rect 11873 15206 11903 15258
rect 11903 15206 11915 15258
rect 11915 15206 11929 15258
rect 11953 15206 11967 15258
rect 11967 15206 11979 15258
rect 11979 15206 12009 15258
rect 12033 15206 12043 15258
rect 12043 15206 12089 15258
rect 11793 15204 11849 15206
rect 11873 15204 11929 15206
rect 11953 15204 12009 15206
rect 12033 15204 12089 15206
rect 11793 14170 11849 14172
rect 11873 14170 11929 14172
rect 11953 14170 12009 14172
rect 12033 14170 12089 14172
rect 11793 14118 11839 14170
rect 11839 14118 11849 14170
rect 11873 14118 11903 14170
rect 11903 14118 11915 14170
rect 11915 14118 11929 14170
rect 11953 14118 11967 14170
rect 11967 14118 11979 14170
rect 11979 14118 12009 14170
rect 12033 14118 12043 14170
rect 12043 14118 12089 14170
rect 11793 14116 11849 14118
rect 11873 14116 11929 14118
rect 11953 14116 12009 14118
rect 12033 14116 12089 14118
rect 15864 17434 15920 17436
rect 15944 17434 16000 17436
rect 16024 17434 16080 17436
rect 16104 17434 16160 17436
rect 15864 17382 15910 17434
rect 15910 17382 15920 17434
rect 15944 17382 15974 17434
rect 15974 17382 15986 17434
rect 15986 17382 16000 17434
rect 16024 17382 16038 17434
rect 16038 17382 16050 17434
rect 16050 17382 16080 17434
rect 16104 17382 16114 17434
rect 16114 17382 16160 17434
rect 15864 17380 15920 17382
rect 15944 17380 16000 17382
rect 16024 17380 16080 17382
rect 16104 17380 16160 17382
rect 15204 16890 15260 16892
rect 15284 16890 15340 16892
rect 15364 16890 15420 16892
rect 15444 16890 15500 16892
rect 15204 16838 15250 16890
rect 15250 16838 15260 16890
rect 15284 16838 15314 16890
rect 15314 16838 15326 16890
rect 15326 16838 15340 16890
rect 15364 16838 15378 16890
rect 15378 16838 15390 16890
rect 15390 16838 15420 16890
rect 15444 16838 15454 16890
rect 15454 16838 15500 16890
rect 15204 16836 15260 16838
rect 15284 16836 15340 16838
rect 15364 16836 15420 16838
rect 15444 16836 15500 16838
rect 15864 16346 15920 16348
rect 15944 16346 16000 16348
rect 16024 16346 16080 16348
rect 16104 16346 16160 16348
rect 15864 16294 15910 16346
rect 15910 16294 15920 16346
rect 15944 16294 15974 16346
rect 15974 16294 15986 16346
rect 15986 16294 16000 16346
rect 16024 16294 16038 16346
rect 16038 16294 16050 16346
rect 16050 16294 16080 16346
rect 16104 16294 16114 16346
rect 16114 16294 16160 16346
rect 15864 16292 15920 16294
rect 15944 16292 16000 16294
rect 16024 16292 16080 16294
rect 16104 16292 16160 16294
rect 15204 15802 15260 15804
rect 15284 15802 15340 15804
rect 15364 15802 15420 15804
rect 15444 15802 15500 15804
rect 15204 15750 15250 15802
rect 15250 15750 15260 15802
rect 15284 15750 15314 15802
rect 15314 15750 15326 15802
rect 15326 15750 15340 15802
rect 15364 15750 15378 15802
rect 15378 15750 15390 15802
rect 15390 15750 15420 15802
rect 15444 15750 15454 15802
rect 15454 15750 15500 15802
rect 15204 15748 15260 15750
rect 15284 15748 15340 15750
rect 15364 15748 15420 15750
rect 15444 15748 15500 15750
rect 11793 13082 11849 13084
rect 11873 13082 11929 13084
rect 11953 13082 12009 13084
rect 12033 13082 12089 13084
rect 11793 13030 11839 13082
rect 11839 13030 11849 13082
rect 11873 13030 11903 13082
rect 11903 13030 11915 13082
rect 11915 13030 11929 13082
rect 11953 13030 11967 13082
rect 11967 13030 11979 13082
rect 11979 13030 12009 13082
rect 12033 13030 12043 13082
rect 12043 13030 12089 13082
rect 11793 13028 11849 13030
rect 11873 13028 11929 13030
rect 11953 13028 12009 13030
rect 12033 13028 12089 13030
rect 15864 15258 15920 15260
rect 15944 15258 16000 15260
rect 16024 15258 16080 15260
rect 16104 15258 16160 15260
rect 15864 15206 15910 15258
rect 15910 15206 15920 15258
rect 15944 15206 15974 15258
rect 15974 15206 15986 15258
rect 15986 15206 16000 15258
rect 16024 15206 16038 15258
rect 16038 15206 16050 15258
rect 16050 15206 16080 15258
rect 16104 15206 16114 15258
rect 16114 15206 16160 15258
rect 15864 15204 15920 15206
rect 15944 15204 16000 15206
rect 16024 15204 16080 15206
rect 16104 15204 16160 15206
rect 15204 14714 15260 14716
rect 15284 14714 15340 14716
rect 15364 14714 15420 14716
rect 15444 14714 15500 14716
rect 15204 14662 15250 14714
rect 15250 14662 15260 14714
rect 15284 14662 15314 14714
rect 15314 14662 15326 14714
rect 15326 14662 15340 14714
rect 15364 14662 15378 14714
rect 15378 14662 15390 14714
rect 15390 14662 15420 14714
rect 15444 14662 15454 14714
rect 15454 14662 15500 14714
rect 15204 14660 15260 14662
rect 15284 14660 15340 14662
rect 15364 14660 15420 14662
rect 15444 14660 15500 14662
rect 15864 14170 15920 14172
rect 15944 14170 16000 14172
rect 16024 14170 16080 14172
rect 16104 14170 16160 14172
rect 15864 14118 15910 14170
rect 15910 14118 15920 14170
rect 15944 14118 15974 14170
rect 15974 14118 15986 14170
rect 15986 14118 16000 14170
rect 16024 14118 16038 14170
rect 16038 14118 16050 14170
rect 16050 14118 16080 14170
rect 16104 14118 16114 14170
rect 16114 14118 16160 14170
rect 15864 14116 15920 14118
rect 15944 14116 16000 14118
rect 16024 14116 16080 14118
rect 16104 14116 16160 14118
rect 16854 15000 16910 15056
rect 17038 14320 17094 14376
rect 7722 10906 7778 10908
rect 7802 10906 7858 10908
rect 7882 10906 7938 10908
rect 7962 10906 8018 10908
rect 7722 10854 7768 10906
rect 7768 10854 7778 10906
rect 7802 10854 7832 10906
rect 7832 10854 7844 10906
rect 7844 10854 7858 10906
rect 7882 10854 7896 10906
rect 7896 10854 7908 10906
rect 7908 10854 7938 10906
rect 7962 10854 7972 10906
rect 7972 10854 8018 10906
rect 7722 10852 7778 10854
rect 7802 10852 7858 10854
rect 7882 10852 7938 10854
rect 7962 10852 8018 10854
rect 3651 8730 3707 8732
rect 3731 8730 3787 8732
rect 3811 8730 3867 8732
rect 3891 8730 3947 8732
rect 3651 8678 3697 8730
rect 3697 8678 3707 8730
rect 3731 8678 3761 8730
rect 3761 8678 3773 8730
rect 3773 8678 3787 8730
rect 3811 8678 3825 8730
rect 3825 8678 3837 8730
rect 3837 8678 3867 8730
rect 3891 8678 3901 8730
rect 3901 8678 3947 8730
rect 3651 8676 3707 8678
rect 3731 8676 3787 8678
rect 3811 8676 3867 8678
rect 3891 8676 3947 8678
rect 2991 8186 3047 8188
rect 3071 8186 3127 8188
rect 3151 8186 3207 8188
rect 3231 8186 3287 8188
rect 2991 8134 3037 8186
rect 3037 8134 3047 8186
rect 3071 8134 3101 8186
rect 3101 8134 3113 8186
rect 3113 8134 3127 8186
rect 3151 8134 3165 8186
rect 3165 8134 3177 8186
rect 3177 8134 3207 8186
rect 3231 8134 3241 8186
rect 3241 8134 3287 8186
rect 2991 8132 3047 8134
rect 3071 8132 3127 8134
rect 3151 8132 3207 8134
rect 3231 8132 3287 8134
rect 2991 7098 3047 7100
rect 3071 7098 3127 7100
rect 3151 7098 3207 7100
rect 3231 7098 3287 7100
rect 2991 7046 3037 7098
rect 3037 7046 3047 7098
rect 3071 7046 3101 7098
rect 3101 7046 3113 7098
rect 3113 7046 3127 7098
rect 3151 7046 3165 7098
rect 3165 7046 3177 7098
rect 3177 7046 3207 7098
rect 3231 7046 3241 7098
rect 3241 7046 3287 7098
rect 2991 7044 3047 7046
rect 3071 7044 3127 7046
rect 3151 7044 3207 7046
rect 3231 7044 3287 7046
rect 3651 7642 3707 7644
rect 3731 7642 3787 7644
rect 3811 7642 3867 7644
rect 3891 7642 3947 7644
rect 3651 7590 3697 7642
rect 3697 7590 3707 7642
rect 3731 7590 3761 7642
rect 3761 7590 3773 7642
rect 3773 7590 3787 7642
rect 3811 7590 3825 7642
rect 3825 7590 3837 7642
rect 3837 7590 3867 7642
rect 3891 7590 3901 7642
rect 3901 7590 3947 7642
rect 3651 7588 3707 7590
rect 3731 7588 3787 7590
rect 3811 7588 3867 7590
rect 3891 7588 3947 7590
rect 4066 6840 4122 6896
rect 2991 6010 3047 6012
rect 3071 6010 3127 6012
rect 3151 6010 3207 6012
rect 3231 6010 3287 6012
rect 2991 5958 3037 6010
rect 3037 5958 3047 6010
rect 3071 5958 3101 6010
rect 3101 5958 3113 6010
rect 3113 5958 3127 6010
rect 3151 5958 3165 6010
rect 3165 5958 3177 6010
rect 3177 5958 3207 6010
rect 3231 5958 3241 6010
rect 3241 5958 3287 6010
rect 2991 5956 3047 5958
rect 3071 5956 3127 5958
rect 3151 5956 3207 5958
rect 3231 5956 3287 5958
rect 3651 6554 3707 6556
rect 3731 6554 3787 6556
rect 3811 6554 3867 6556
rect 3891 6554 3947 6556
rect 3651 6502 3697 6554
rect 3697 6502 3707 6554
rect 3731 6502 3761 6554
rect 3761 6502 3773 6554
rect 3773 6502 3787 6554
rect 3811 6502 3825 6554
rect 3825 6502 3837 6554
rect 3837 6502 3867 6554
rect 3891 6502 3901 6554
rect 3901 6502 3947 6554
rect 3651 6500 3707 6502
rect 3731 6500 3787 6502
rect 3811 6500 3867 6502
rect 3891 6500 3947 6502
rect 3651 5466 3707 5468
rect 3731 5466 3787 5468
rect 3811 5466 3867 5468
rect 3891 5466 3947 5468
rect 3651 5414 3697 5466
rect 3697 5414 3707 5466
rect 3731 5414 3761 5466
rect 3761 5414 3773 5466
rect 3773 5414 3787 5466
rect 3811 5414 3825 5466
rect 3825 5414 3837 5466
rect 3837 5414 3867 5466
rect 3891 5414 3901 5466
rect 3901 5414 3947 5466
rect 3651 5412 3707 5414
rect 3731 5412 3787 5414
rect 3811 5412 3867 5414
rect 3891 5412 3947 5414
rect 7062 10362 7118 10364
rect 7142 10362 7198 10364
rect 7222 10362 7278 10364
rect 7302 10362 7358 10364
rect 7062 10310 7108 10362
rect 7108 10310 7118 10362
rect 7142 10310 7172 10362
rect 7172 10310 7184 10362
rect 7184 10310 7198 10362
rect 7222 10310 7236 10362
rect 7236 10310 7248 10362
rect 7248 10310 7278 10362
rect 7302 10310 7312 10362
rect 7312 10310 7358 10362
rect 7062 10308 7118 10310
rect 7142 10308 7198 10310
rect 7222 10308 7278 10310
rect 7302 10308 7358 10310
rect 7062 9274 7118 9276
rect 7142 9274 7198 9276
rect 7222 9274 7278 9276
rect 7302 9274 7358 9276
rect 7062 9222 7108 9274
rect 7108 9222 7118 9274
rect 7142 9222 7172 9274
rect 7172 9222 7184 9274
rect 7184 9222 7198 9274
rect 7222 9222 7236 9274
rect 7236 9222 7248 9274
rect 7248 9222 7278 9274
rect 7302 9222 7312 9274
rect 7312 9222 7358 9274
rect 7062 9220 7118 9222
rect 7142 9220 7198 9222
rect 7222 9220 7278 9222
rect 7302 9220 7358 9222
rect 7062 8186 7118 8188
rect 7142 8186 7198 8188
rect 7222 8186 7278 8188
rect 7302 8186 7358 8188
rect 7062 8134 7108 8186
rect 7108 8134 7118 8186
rect 7142 8134 7172 8186
rect 7172 8134 7184 8186
rect 7184 8134 7198 8186
rect 7222 8134 7236 8186
rect 7236 8134 7248 8186
rect 7248 8134 7278 8186
rect 7302 8134 7312 8186
rect 7312 8134 7358 8186
rect 7062 8132 7118 8134
rect 7142 8132 7198 8134
rect 7222 8132 7278 8134
rect 7302 8132 7358 8134
rect 7722 9818 7778 9820
rect 7802 9818 7858 9820
rect 7882 9818 7938 9820
rect 7962 9818 8018 9820
rect 7722 9766 7768 9818
rect 7768 9766 7778 9818
rect 7802 9766 7832 9818
rect 7832 9766 7844 9818
rect 7844 9766 7858 9818
rect 7882 9766 7896 9818
rect 7896 9766 7908 9818
rect 7908 9766 7938 9818
rect 7962 9766 7972 9818
rect 7972 9766 8018 9818
rect 7722 9764 7778 9766
rect 7802 9764 7858 9766
rect 7882 9764 7938 9766
rect 7962 9764 8018 9766
rect 7722 8730 7778 8732
rect 7802 8730 7858 8732
rect 7882 8730 7938 8732
rect 7962 8730 8018 8732
rect 7722 8678 7768 8730
rect 7768 8678 7778 8730
rect 7802 8678 7832 8730
rect 7832 8678 7844 8730
rect 7844 8678 7858 8730
rect 7882 8678 7896 8730
rect 7896 8678 7908 8730
rect 7908 8678 7938 8730
rect 7962 8678 7972 8730
rect 7972 8678 8018 8730
rect 7722 8676 7778 8678
rect 7802 8676 7858 8678
rect 7882 8676 7938 8678
rect 7962 8676 8018 8678
rect 11133 12538 11189 12540
rect 11213 12538 11269 12540
rect 11293 12538 11349 12540
rect 11373 12538 11429 12540
rect 11133 12486 11179 12538
rect 11179 12486 11189 12538
rect 11213 12486 11243 12538
rect 11243 12486 11255 12538
rect 11255 12486 11269 12538
rect 11293 12486 11307 12538
rect 11307 12486 11319 12538
rect 11319 12486 11349 12538
rect 11373 12486 11383 12538
rect 11383 12486 11429 12538
rect 11133 12484 11189 12486
rect 11213 12484 11269 12486
rect 11293 12484 11349 12486
rect 11373 12484 11429 12486
rect 11793 11994 11849 11996
rect 11873 11994 11929 11996
rect 11953 11994 12009 11996
rect 12033 11994 12089 11996
rect 11793 11942 11839 11994
rect 11839 11942 11849 11994
rect 11873 11942 11903 11994
rect 11903 11942 11915 11994
rect 11915 11942 11929 11994
rect 11953 11942 11967 11994
rect 11967 11942 11979 11994
rect 11979 11942 12009 11994
rect 12033 11942 12043 11994
rect 12043 11942 12089 11994
rect 11793 11940 11849 11942
rect 11873 11940 11929 11942
rect 11953 11940 12009 11942
rect 12033 11940 12089 11942
rect 15204 13626 15260 13628
rect 15284 13626 15340 13628
rect 15364 13626 15420 13628
rect 15444 13626 15500 13628
rect 15204 13574 15250 13626
rect 15250 13574 15260 13626
rect 15284 13574 15314 13626
rect 15314 13574 15326 13626
rect 15326 13574 15340 13626
rect 15364 13574 15378 13626
rect 15378 13574 15390 13626
rect 15390 13574 15420 13626
rect 15444 13574 15454 13626
rect 15454 13574 15500 13626
rect 15204 13572 15260 13574
rect 15284 13572 15340 13574
rect 15364 13572 15420 13574
rect 15444 13572 15500 13574
rect 15864 13082 15920 13084
rect 15944 13082 16000 13084
rect 16024 13082 16080 13084
rect 16104 13082 16160 13084
rect 15864 13030 15910 13082
rect 15910 13030 15920 13082
rect 15944 13030 15974 13082
rect 15974 13030 15986 13082
rect 15986 13030 16000 13082
rect 16024 13030 16038 13082
rect 16038 13030 16050 13082
rect 16050 13030 16080 13082
rect 16104 13030 16114 13082
rect 16114 13030 16160 13082
rect 15864 13028 15920 13030
rect 15944 13028 16000 13030
rect 16024 13028 16080 13030
rect 16104 13028 16160 13030
rect 11133 11450 11189 11452
rect 11213 11450 11269 11452
rect 11293 11450 11349 11452
rect 11373 11450 11429 11452
rect 11133 11398 11179 11450
rect 11179 11398 11189 11450
rect 11213 11398 11243 11450
rect 11243 11398 11255 11450
rect 11255 11398 11269 11450
rect 11293 11398 11307 11450
rect 11307 11398 11319 11450
rect 11319 11398 11349 11450
rect 11373 11398 11383 11450
rect 11383 11398 11429 11450
rect 11133 11396 11189 11398
rect 11213 11396 11269 11398
rect 11293 11396 11349 11398
rect 11373 11396 11429 11398
rect 11793 10906 11849 10908
rect 11873 10906 11929 10908
rect 11953 10906 12009 10908
rect 12033 10906 12089 10908
rect 11793 10854 11839 10906
rect 11839 10854 11849 10906
rect 11873 10854 11903 10906
rect 11903 10854 11915 10906
rect 11915 10854 11929 10906
rect 11953 10854 11967 10906
rect 11967 10854 11979 10906
rect 11979 10854 12009 10906
rect 12033 10854 12043 10906
rect 12043 10854 12089 10906
rect 11793 10852 11849 10854
rect 11873 10852 11929 10854
rect 11953 10852 12009 10854
rect 12033 10852 12089 10854
rect 15204 12538 15260 12540
rect 15284 12538 15340 12540
rect 15364 12538 15420 12540
rect 15444 12538 15500 12540
rect 15204 12486 15250 12538
rect 15250 12486 15260 12538
rect 15284 12486 15314 12538
rect 15314 12486 15326 12538
rect 15326 12486 15340 12538
rect 15364 12486 15378 12538
rect 15378 12486 15390 12538
rect 15390 12486 15420 12538
rect 15444 12486 15454 12538
rect 15454 12486 15500 12538
rect 15204 12484 15260 12486
rect 15284 12484 15340 12486
rect 15364 12484 15420 12486
rect 15444 12484 15500 12486
rect 17038 12960 17094 13016
rect 15864 11994 15920 11996
rect 15944 11994 16000 11996
rect 16024 11994 16080 11996
rect 16104 11994 16160 11996
rect 15864 11942 15910 11994
rect 15910 11942 15920 11994
rect 15944 11942 15974 11994
rect 15974 11942 15986 11994
rect 15986 11942 16000 11994
rect 16024 11942 16038 11994
rect 16038 11942 16050 11994
rect 16050 11942 16080 11994
rect 16104 11942 16114 11994
rect 16114 11942 16160 11994
rect 15864 11940 15920 11942
rect 15944 11940 16000 11942
rect 16024 11940 16080 11942
rect 16104 11940 16160 11942
rect 15204 11450 15260 11452
rect 15284 11450 15340 11452
rect 15364 11450 15420 11452
rect 15444 11450 15500 11452
rect 15204 11398 15250 11450
rect 15250 11398 15260 11450
rect 15284 11398 15314 11450
rect 15314 11398 15326 11450
rect 15326 11398 15340 11450
rect 15364 11398 15378 11450
rect 15378 11398 15390 11450
rect 15390 11398 15420 11450
rect 15444 11398 15454 11450
rect 15454 11398 15500 11450
rect 15204 11396 15260 11398
rect 15284 11396 15340 11398
rect 15364 11396 15420 11398
rect 15444 11396 15500 11398
rect 11133 10362 11189 10364
rect 11213 10362 11269 10364
rect 11293 10362 11349 10364
rect 11373 10362 11429 10364
rect 11133 10310 11179 10362
rect 11179 10310 11189 10362
rect 11213 10310 11243 10362
rect 11243 10310 11255 10362
rect 11255 10310 11269 10362
rect 11293 10310 11307 10362
rect 11307 10310 11319 10362
rect 11319 10310 11349 10362
rect 11373 10310 11383 10362
rect 11383 10310 11429 10362
rect 11133 10308 11189 10310
rect 11213 10308 11269 10310
rect 11293 10308 11349 10310
rect 11373 10308 11429 10310
rect 7062 7098 7118 7100
rect 7142 7098 7198 7100
rect 7222 7098 7278 7100
rect 7302 7098 7358 7100
rect 7062 7046 7108 7098
rect 7108 7046 7118 7098
rect 7142 7046 7172 7098
rect 7172 7046 7184 7098
rect 7184 7046 7198 7098
rect 7222 7046 7236 7098
rect 7236 7046 7248 7098
rect 7248 7046 7278 7098
rect 7302 7046 7312 7098
rect 7312 7046 7358 7098
rect 7062 7044 7118 7046
rect 7142 7044 7198 7046
rect 7222 7044 7278 7046
rect 7302 7044 7358 7046
rect 7062 6010 7118 6012
rect 7142 6010 7198 6012
rect 7222 6010 7278 6012
rect 7302 6010 7358 6012
rect 7062 5958 7108 6010
rect 7108 5958 7118 6010
rect 7142 5958 7172 6010
rect 7172 5958 7184 6010
rect 7184 5958 7198 6010
rect 7222 5958 7236 6010
rect 7236 5958 7248 6010
rect 7248 5958 7278 6010
rect 7302 5958 7312 6010
rect 7312 5958 7358 6010
rect 7062 5956 7118 5958
rect 7142 5956 7198 5958
rect 7222 5956 7278 5958
rect 7302 5956 7358 5958
rect 2991 4922 3047 4924
rect 3071 4922 3127 4924
rect 3151 4922 3207 4924
rect 3231 4922 3287 4924
rect 2991 4870 3037 4922
rect 3037 4870 3047 4922
rect 3071 4870 3101 4922
rect 3101 4870 3113 4922
rect 3113 4870 3127 4922
rect 3151 4870 3165 4922
rect 3165 4870 3177 4922
rect 3177 4870 3207 4922
rect 3231 4870 3241 4922
rect 3241 4870 3287 4922
rect 2991 4868 3047 4870
rect 3071 4868 3127 4870
rect 3151 4868 3207 4870
rect 3231 4868 3287 4870
rect 3651 4378 3707 4380
rect 3731 4378 3787 4380
rect 3811 4378 3867 4380
rect 3891 4378 3947 4380
rect 3651 4326 3697 4378
rect 3697 4326 3707 4378
rect 3731 4326 3761 4378
rect 3761 4326 3773 4378
rect 3773 4326 3787 4378
rect 3811 4326 3825 4378
rect 3825 4326 3837 4378
rect 3837 4326 3867 4378
rect 3891 4326 3901 4378
rect 3901 4326 3947 4378
rect 3651 4324 3707 4326
rect 3731 4324 3787 4326
rect 3811 4324 3867 4326
rect 3891 4324 3947 4326
rect 2991 3834 3047 3836
rect 3071 3834 3127 3836
rect 3151 3834 3207 3836
rect 3231 3834 3287 3836
rect 2991 3782 3037 3834
rect 3037 3782 3047 3834
rect 3071 3782 3101 3834
rect 3101 3782 3113 3834
rect 3113 3782 3127 3834
rect 3151 3782 3165 3834
rect 3165 3782 3177 3834
rect 3177 3782 3207 3834
rect 3231 3782 3241 3834
rect 3241 3782 3287 3834
rect 2991 3780 3047 3782
rect 3071 3780 3127 3782
rect 3151 3780 3207 3782
rect 3231 3780 3287 3782
rect 3651 3290 3707 3292
rect 3731 3290 3787 3292
rect 3811 3290 3867 3292
rect 3891 3290 3947 3292
rect 3651 3238 3697 3290
rect 3697 3238 3707 3290
rect 3731 3238 3761 3290
rect 3761 3238 3773 3290
rect 3773 3238 3787 3290
rect 3811 3238 3825 3290
rect 3825 3238 3837 3290
rect 3837 3238 3867 3290
rect 3891 3238 3901 3290
rect 3901 3238 3947 3290
rect 3651 3236 3707 3238
rect 3731 3236 3787 3238
rect 3811 3236 3867 3238
rect 3891 3236 3947 3238
rect 2991 2746 3047 2748
rect 3071 2746 3127 2748
rect 3151 2746 3207 2748
rect 3231 2746 3287 2748
rect 2991 2694 3037 2746
rect 3037 2694 3047 2746
rect 3071 2694 3101 2746
rect 3101 2694 3113 2746
rect 3113 2694 3127 2746
rect 3151 2694 3165 2746
rect 3165 2694 3177 2746
rect 3177 2694 3207 2746
rect 3231 2694 3241 2746
rect 3241 2694 3287 2746
rect 2991 2692 3047 2694
rect 3071 2692 3127 2694
rect 3151 2692 3207 2694
rect 3231 2692 3287 2694
rect 7722 7642 7778 7644
rect 7802 7642 7858 7644
rect 7882 7642 7938 7644
rect 7962 7642 8018 7644
rect 7722 7590 7768 7642
rect 7768 7590 7778 7642
rect 7802 7590 7832 7642
rect 7832 7590 7844 7642
rect 7844 7590 7858 7642
rect 7882 7590 7896 7642
rect 7896 7590 7908 7642
rect 7908 7590 7938 7642
rect 7962 7590 7972 7642
rect 7972 7590 8018 7642
rect 7722 7588 7778 7590
rect 7802 7588 7858 7590
rect 7882 7588 7938 7590
rect 7962 7588 8018 7590
rect 11793 9818 11849 9820
rect 11873 9818 11929 9820
rect 11953 9818 12009 9820
rect 12033 9818 12089 9820
rect 11793 9766 11839 9818
rect 11839 9766 11849 9818
rect 11873 9766 11903 9818
rect 11903 9766 11915 9818
rect 11915 9766 11929 9818
rect 11953 9766 11967 9818
rect 11967 9766 11979 9818
rect 11979 9766 12009 9818
rect 12033 9766 12043 9818
rect 12043 9766 12089 9818
rect 11793 9764 11849 9766
rect 11873 9764 11929 9766
rect 11953 9764 12009 9766
rect 12033 9764 12089 9766
rect 11133 9274 11189 9276
rect 11213 9274 11269 9276
rect 11293 9274 11349 9276
rect 11373 9274 11429 9276
rect 11133 9222 11179 9274
rect 11179 9222 11189 9274
rect 11213 9222 11243 9274
rect 11243 9222 11255 9274
rect 11255 9222 11269 9274
rect 11293 9222 11307 9274
rect 11307 9222 11319 9274
rect 11319 9222 11349 9274
rect 11373 9222 11383 9274
rect 11383 9222 11429 9274
rect 11133 9220 11189 9222
rect 11213 9220 11269 9222
rect 11293 9220 11349 9222
rect 11373 9220 11429 9222
rect 11793 8730 11849 8732
rect 11873 8730 11929 8732
rect 11953 8730 12009 8732
rect 12033 8730 12089 8732
rect 11793 8678 11839 8730
rect 11839 8678 11849 8730
rect 11873 8678 11903 8730
rect 11903 8678 11915 8730
rect 11915 8678 11929 8730
rect 11953 8678 11967 8730
rect 11967 8678 11979 8730
rect 11979 8678 12009 8730
rect 12033 8678 12043 8730
rect 12043 8678 12089 8730
rect 11793 8676 11849 8678
rect 11873 8676 11929 8678
rect 11953 8676 12009 8678
rect 12033 8676 12089 8678
rect 7722 6554 7778 6556
rect 7802 6554 7858 6556
rect 7882 6554 7938 6556
rect 7962 6554 8018 6556
rect 7722 6502 7768 6554
rect 7768 6502 7778 6554
rect 7802 6502 7832 6554
rect 7832 6502 7844 6554
rect 7844 6502 7858 6554
rect 7882 6502 7896 6554
rect 7896 6502 7908 6554
rect 7908 6502 7938 6554
rect 7962 6502 7972 6554
rect 7972 6502 8018 6554
rect 7722 6500 7778 6502
rect 7802 6500 7858 6502
rect 7882 6500 7938 6502
rect 7962 6500 8018 6502
rect 7722 5466 7778 5468
rect 7802 5466 7858 5468
rect 7882 5466 7938 5468
rect 7962 5466 8018 5468
rect 7722 5414 7768 5466
rect 7768 5414 7778 5466
rect 7802 5414 7832 5466
rect 7832 5414 7844 5466
rect 7844 5414 7858 5466
rect 7882 5414 7896 5466
rect 7896 5414 7908 5466
rect 7908 5414 7938 5466
rect 7962 5414 7972 5466
rect 7972 5414 8018 5466
rect 7722 5412 7778 5414
rect 7802 5412 7858 5414
rect 7882 5412 7938 5414
rect 7962 5412 8018 5414
rect 7062 4922 7118 4924
rect 7142 4922 7198 4924
rect 7222 4922 7278 4924
rect 7302 4922 7358 4924
rect 7062 4870 7108 4922
rect 7108 4870 7118 4922
rect 7142 4870 7172 4922
rect 7172 4870 7184 4922
rect 7184 4870 7198 4922
rect 7222 4870 7236 4922
rect 7236 4870 7248 4922
rect 7248 4870 7278 4922
rect 7302 4870 7312 4922
rect 7312 4870 7358 4922
rect 7062 4868 7118 4870
rect 7142 4868 7198 4870
rect 7222 4868 7278 4870
rect 7302 4868 7358 4870
rect 7722 4378 7778 4380
rect 7802 4378 7858 4380
rect 7882 4378 7938 4380
rect 7962 4378 8018 4380
rect 7722 4326 7768 4378
rect 7768 4326 7778 4378
rect 7802 4326 7832 4378
rect 7832 4326 7844 4378
rect 7844 4326 7858 4378
rect 7882 4326 7896 4378
rect 7896 4326 7908 4378
rect 7908 4326 7938 4378
rect 7962 4326 7972 4378
rect 7972 4326 8018 4378
rect 7722 4324 7778 4326
rect 7802 4324 7858 4326
rect 7882 4324 7938 4326
rect 7962 4324 8018 4326
rect 7062 3834 7118 3836
rect 7142 3834 7198 3836
rect 7222 3834 7278 3836
rect 7302 3834 7358 3836
rect 7062 3782 7108 3834
rect 7108 3782 7118 3834
rect 7142 3782 7172 3834
rect 7172 3782 7184 3834
rect 7184 3782 7198 3834
rect 7222 3782 7236 3834
rect 7236 3782 7248 3834
rect 7248 3782 7278 3834
rect 7302 3782 7312 3834
rect 7312 3782 7358 3834
rect 7062 3780 7118 3782
rect 7142 3780 7198 3782
rect 7222 3780 7278 3782
rect 7302 3780 7358 3782
rect 7722 3290 7778 3292
rect 7802 3290 7858 3292
rect 7882 3290 7938 3292
rect 7962 3290 8018 3292
rect 7722 3238 7768 3290
rect 7768 3238 7778 3290
rect 7802 3238 7832 3290
rect 7832 3238 7844 3290
rect 7844 3238 7858 3290
rect 7882 3238 7896 3290
rect 7896 3238 7908 3290
rect 7908 3238 7938 3290
rect 7962 3238 7972 3290
rect 7972 3238 8018 3290
rect 7722 3236 7778 3238
rect 7802 3236 7858 3238
rect 7882 3236 7938 3238
rect 7962 3236 8018 3238
rect 7062 2746 7118 2748
rect 7142 2746 7198 2748
rect 7222 2746 7278 2748
rect 7302 2746 7358 2748
rect 7062 2694 7108 2746
rect 7108 2694 7118 2746
rect 7142 2694 7172 2746
rect 7172 2694 7184 2746
rect 7184 2694 7198 2746
rect 7222 2694 7236 2746
rect 7236 2694 7248 2746
rect 7248 2694 7278 2746
rect 7302 2694 7312 2746
rect 7312 2694 7358 2746
rect 7062 2692 7118 2694
rect 7142 2692 7198 2694
rect 7222 2692 7278 2694
rect 7302 2692 7358 2694
rect 11133 8186 11189 8188
rect 11213 8186 11269 8188
rect 11293 8186 11349 8188
rect 11373 8186 11429 8188
rect 11133 8134 11179 8186
rect 11179 8134 11189 8186
rect 11213 8134 11243 8186
rect 11243 8134 11255 8186
rect 11255 8134 11269 8186
rect 11293 8134 11307 8186
rect 11307 8134 11319 8186
rect 11319 8134 11349 8186
rect 11373 8134 11383 8186
rect 11383 8134 11429 8186
rect 11133 8132 11189 8134
rect 11213 8132 11269 8134
rect 11293 8132 11349 8134
rect 11373 8132 11429 8134
rect 11793 7642 11849 7644
rect 11873 7642 11929 7644
rect 11953 7642 12009 7644
rect 12033 7642 12089 7644
rect 11793 7590 11839 7642
rect 11839 7590 11849 7642
rect 11873 7590 11903 7642
rect 11903 7590 11915 7642
rect 11915 7590 11929 7642
rect 11953 7590 11967 7642
rect 11967 7590 11979 7642
rect 11979 7590 12009 7642
rect 12033 7590 12043 7642
rect 12043 7590 12089 7642
rect 11793 7588 11849 7590
rect 11873 7588 11929 7590
rect 11953 7588 12009 7590
rect 12033 7588 12089 7590
rect 15204 10362 15260 10364
rect 15284 10362 15340 10364
rect 15364 10362 15420 10364
rect 15444 10362 15500 10364
rect 15204 10310 15250 10362
rect 15250 10310 15260 10362
rect 15284 10310 15314 10362
rect 15314 10310 15326 10362
rect 15326 10310 15340 10362
rect 15364 10310 15378 10362
rect 15378 10310 15390 10362
rect 15390 10310 15420 10362
rect 15444 10310 15454 10362
rect 15454 10310 15500 10362
rect 15204 10308 15260 10310
rect 15284 10308 15340 10310
rect 15364 10308 15420 10310
rect 15444 10308 15500 10310
rect 15864 10906 15920 10908
rect 15944 10906 16000 10908
rect 16024 10906 16080 10908
rect 16104 10906 16160 10908
rect 15864 10854 15910 10906
rect 15910 10854 15920 10906
rect 15944 10854 15974 10906
rect 15974 10854 15986 10906
rect 15986 10854 16000 10906
rect 16024 10854 16038 10906
rect 16038 10854 16050 10906
rect 16050 10854 16080 10906
rect 16104 10854 16114 10906
rect 16114 10854 16160 10906
rect 15864 10852 15920 10854
rect 15944 10852 16000 10854
rect 16024 10852 16080 10854
rect 16104 10852 16160 10854
rect 16486 11600 16542 11656
rect 11133 7098 11189 7100
rect 11213 7098 11269 7100
rect 11293 7098 11349 7100
rect 11373 7098 11429 7100
rect 11133 7046 11179 7098
rect 11179 7046 11189 7098
rect 11213 7046 11243 7098
rect 11243 7046 11255 7098
rect 11255 7046 11269 7098
rect 11293 7046 11307 7098
rect 11307 7046 11319 7098
rect 11319 7046 11349 7098
rect 11373 7046 11383 7098
rect 11383 7046 11429 7098
rect 11133 7044 11189 7046
rect 11213 7044 11269 7046
rect 11293 7044 11349 7046
rect 11373 7044 11429 7046
rect 11133 6010 11189 6012
rect 11213 6010 11269 6012
rect 11293 6010 11349 6012
rect 11373 6010 11429 6012
rect 11133 5958 11179 6010
rect 11179 5958 11189 6010
rect 11213 5958 11243 6010
rect 11243 5958 11255 6010
rect 11255 5958 11269 6010
rect 11293 5958 11307 6010
rect 11307 5958 11319 6010
rect 11319 5958 11349 6010
rect 11373 5958 11383 6010
rect 11383 5958 11429 6010
rect 11133 5956 11189 5958
rect 11213 5956 11269 5958
rect 11293 5956 11349 5958
rect 11373 5956 11429 5958
rect 11793 6554 11849 6556
rect 11873 6554 11929 6556
rect 11953 6554 12009 6556
rect 12033 6554 12089 6556
rect 11793 6502 11839 6554
rect 11839 6502 11849 6554
rect 11873 6502 11903 6554
rect 11903 6502 11915 6554
rect 11915 6502 11929 6554
rect 11953 6502 11967 6554
rect 11967 6502 11979 6554
rect 11979 6502 12009 6554
rect 12033 6502 12043 6554
rect 12043 6502 12089 6554
rect 11793 6500 11849 6502
rect 11873 6500 11929 6502
rect 11953 6500 12009 6502
rect 12033 6500 12089 6502
rect 11133 4922 11189 4924
rect 11213 4922 11269 4924
rect 11293 4922 11349 4924
rect 11373 4922 11429 4924
rect 11133 4870 11179 4922
rect 11179 4870 11189 4922
rect 11213 4870 11243 4922
rect 11243 4870 11255 4922
rect 11255 4870 11269 4922
rect 11293 4870 11307 4922
rect 11307 4870 11319 4922
rect 11319 4870 11349 4922
rect 11373 4870 11383 4922
rect 11383 4870 11429 4922
rect 11133 4868 11189 4870
rect 11213 4868 11269 4870
rect 11293 4868 11349 4870
rect 11373 4868 11429 4870
rect 11133 3834 11189 3836
rect 11213 3834 11269 3836
rect 11293 3834 11349 3836
rect 11373 3834 11429 3836
rect 11133 3782 11179 3834
rect 11179 3782 11189 3834
rect 11213 3782 11243 3834
rect 11243 3782 11255 3834
rect 11255 3782 11269 3834
rect 11293 3782 11307 3834
rect 11307 3782 11319 3834
rect 11319 3782 11349 3834
rect 11373 3782 11383 3834
rect 11383 3782 11429 3834
rect 11133 3780 11189 3782
rect 11213 3780 11269 3782
rect 11293 3780 11349 3782
rect 11373 3780 11429 3782
rect 11133 2746 11189 2748
rect 11213 2746 11269 2748
rect 11293 2746 11349 2748
rect 11373 2746 11429 2748
rect 11133 2694 11179 2746
rect 11179 2694 11189 2746
rect 11213 2694 11243 2746
rect 11243 2694 11255 2746
rect 11255 2694 11269 2746
rect 11293 2694 11307 2746
rect 11307 2694 11319 2746
rect 11319 2694 11349 2746
rect 11373 2694 11383 2746
rect 11383 2694 11429 2746
rect 11133 2692 11189 2694
rect 11213 2692 11269 2694
rect 11293 2692 11349 2694
rect 11373 2692 11429 2694
rect 15204 9274 15260 9276
rect 15284 9274 15340 9276
rect 15364 9274 15420 9276
rect 15444 9274 15500 9276
rect 15204 9222 15250 9274
rect 15250 9222 15260 9274
rect 15284 9222 15314 9274
rect 15314 9222 15326 9274
rect 15326 9222 15340 9274
rect 15364 9222 15378 9274
rect 15378 9222 15390 9274
rect 15390 9222 15420 9274
rect 15444 9222 15454 9274
rect 15454 9222 15500 9274
rect 15204 9220 15260 9222
rect 15284 9220 15340 9222
rect 15364 9220 15420 9222
rect 15444 9220 15500 9222
rect 15864 9818 15920 9820
rect 15944 9818 16000 9820
rect 16024 9818 16080 9820
rect 16104 9818 16160 9820
rect 15864 9766 15910 9818
rect 15910 9766 15920 9818
rect 15944 9766 15974 9818
rect 15974 9766 15986 9818
rect 15986 9766 16000 9818
rect 16024 9766 16038 9818
rect 16038 9766 16050 9818
rect 16050 9766 16080 9818
rect 16104 9766 16114 9818
rect 16114 9766 16160 9818
rect 15864 9764 15920 9766
rect 15944 9764 16000 9766
rect 16024 9764 16080 9766
rect 16104 9764 16160 9766
rect 17038 10920 17094 10976
rect 15864 8730 15920 8732
rect 15944 8730 16000 8732
rect 16024 8730 16080 8732
rect 16104 8730 16160 8732
rect 15864 8678 15910 8730
rect 15910 8678 15920 8730
rect 15944 8678 15974 8730
rect 15974 8678 15986 8730
rect 15986 8678 16000 8730
rect 16024 8678 16038 8730
rect 16038 8678 16050 8730
rect 16050 8678 16080 8730
rect 16104 8678 16114 8730
rect 16114 8678 16160 8730
rect 15864 8676 15920 8678
rect 15944 8676 16000 8678
rect 16024 8676 16080 8678
rect 16104 8676 16160 8678
rect 15204 8186 15260 8188
rect 15284 8186 15340 8188
rect 15364 8186 15420 8188
rect 15444 8186 15500 8188
rect 15204 8134 15250 8186
rect 15250 8134 15260 8186
rect 15284 8134 15314 8186
rect 15314 8134 15326 8186
rect 15326 8134 15340 8186
rect 15364 8134 15378 8186
rect 15378 8134 15390 8186
rect 15390 8134 15420 8186
rect 15444 8134 15454 8186
rect 15454 8134 15500 8186
rect 15204 8132 15260 8134
rect 15284 8132 15340 8134
rect 15364 8132 15420 8134
rect 15444 8132 15500 8134
rect 15864 7642 15920 7644
rect 15944 7642 16000 7644
rect 16024 7642 16080 7644
rect 16104 7642 16160 7644
rect 15864 7590 15910 7642
rect 15910 7590 15920 7642
rect 15944 7590 15974 7642
rect 15974 7590 15986 7642
rect 15986 7590 16000 7642
rect 16024 7590 16038 7642
rect 16038 7590 16050 7642
rect 16050 7590 16080 7642
rect 16104 7590 16114 7642
rect 16114 7590 16160 7642
rect 15864 7588 15920 7590
rect 15944 7588 16000 7590
rect 16024 7588 16080 7590
rect 16104 7588 16160 7590
rect 11793 5466 11849 5468
rect 11873 5466 11929 5468
rect 11953 5466 12009 5468
rect 12033 5466 12089 5468
rect 11793 5414 11839 5466
rect 11839 5414 11849 5466
rect 11873 5414 11903 5466
rect 11903 5414 11915 5466
rect 11915 5414 11929 5466
rect 11953 5414 11967 5466
rect 11967 5414 11979 5466
rect 11979 5414 12009 5466
rect 12033 5414 12043 5466
rect 12043 5414 12089 5466
rect 11793 5412 11849 5414
rect 11873 5412 11929 5414
rect 11953 5412 12009 5414
rect 12033 5412 12089 5414
rect 11793 4378 11849 4380
rect 11873 4378 11929 4380
rect 11953 4378 12009 4380
rect 12033 4378 12089 4380
rect 11793 4326 11839 4378
rect 11839 4326 11849 4378
rect 11873 4326 11903 4378
rect 11903 4326 11915 4378
rect 11915 4326 11929 4378
rect 11953 4326 11967 4378
rect 11967 4326 11979 4378
rect 11979 4326 12009 4378
rect 12033 4326 12043 4378
rect 12043 4326 12089 4378
rect 11793 4324 11849 4326
rect 11873 4324 11929 4326
rect 11953 4324 12009 4326
rect 12033 4324 12089 4326
rect 11793 3290 11849 3292
rect 11873 3290 11929 3292
rect 11953 3290 12009 3292
rect 12033 3290 12089 3292
rect 11793 3238 11839 3290
rect 11839 3238 11849 3290
rect 11873 3238 11903 3290
rect 11903 3238 11915 3290
rect 11915 3238 11929 3290
rect 11953 3238 11967 3290
rect 11967 3238 11979 3290
rect 11979 3238 12009 3290
rect 12033 3238 12043 3290
rect 12043 3238 12089 3290
rect 11793 3236 11849 3238
rect 11873 3236 11929 3238
rect 11953 3236 12009 3238
rect 12033 3236 12089 3238
rect 15204 7098 15260 7100
rect 15284 7098 15340 7100
rect 15364 7098 15420 7100
rect 15444 7098 15500 7100
rect 15204 7046 15250 7098
rect 15250 7046 15260 7098
rect 15284 7046 15314 7098
rect 15314 7046 15326 7098
rect 15326 7046 15340 7098
rect 15364 7046 15378 7098
rect 15378 7046 15390 7098
rect 15390 7046 15420 7098
rect 15444 7046 15454 7098
rect 15454 7046 15500 7098
rect 15204 7044 15260 7046
rect 15284 7044 15340 7046
rect 15364 7044 15420 7046
rect 15444 7044 15500 7046
rect 15204 6010 15260 6012
rect 15284 6010 15340 6012
rect 15364 6010 15420 6012
rect 15444 6010 15500 6012
rect 15204 5958 15250 6010
rect 15250 5958 15260 6010
rect 15284 5958 15314 6010
rect 15314 5958 15326 6010
rect 15326 5958 15340 6010
rect 15364 5958 15378 6010
rect 15378 5958 15390 6010
rect 15390 5958 15420 6010
rect 15444 5958 15454 6010
rect 15454 5958 15500 6010
rect 15204 5956 15260 5958
rect 15284 5956 15340 5958
rect 15364 5956 15420 5958
rect 15444 5956 15500 5958
rect 15864 6554 15920 6556
rect 15944 6554 16000 6556
rect 16024 6554 16080 6556
rect 16104 6554 16160 6556
rect 15864 6502 15910 6554
rect 15910 6502 15920 6554
rect 15944 6502 15974 6554
rect 15974 6502 15986 6554
rect 15986 6502 16000 6554
rect 16024 6502 16038 6554
rect 16038 6502 16050 6554
rect 16050 6502 16080 6554
rect 16104 6502 16114 6554
rect 16114 6502 16160 6554
rect 15864 6500 15920 6502
rect 15944 6500 16000 6502
rect 16024 6500 16080 6502
rect 16104 6500 16160 6502
rect 15864 5466 15920 5468
rect 15944 5466 16000 5468
rect 16024 5466 16080 5468
rect 16104 5466 16160 5468
rect 15864 5414 15910 5466
rect 15910 5414 15920 5466
rect 15944 5414 15974 5466
rect 15974 5414 15986 5466
rect 15986 5414 16000 5466
rect 16024 5414 16038 5466
rect 16038 5414 16050 5466
rect 16050 5414 16080 5466
rect 16104 5414 16114 5466
rect 16114 5414 16160 5466
rect 15864 5412 15920 5414
rect 15944 5412 16000 5414
rect 16024 5412 16080 5414
rect 16104 5412 16160 5414
rect 15204 4922 15260 4924
rect 15284 4922 15340 4924
rect 15364 4922 15420 4924
rect 15444 4922 15500 4924
rect 15204 4870 15250 4922
rect 15250 4870 15260 4922
rect 15284 4870 15314 4922
rect 15314 4870 15326 4922
rect 15326 4870 15340 4922
rect 15364 4870 15378 4922
rect 15378 4870 15390 4922
rect 15390 4870 15420 4922
rect 15444 4870 15454 4922
rect 15454 4870 15500 4922
rect 15204 4868 15260 4870
rect 15284 4868 15340 4870
rect 15364 4868 15420 4870
rect 15444 4868 15500 4870
rect 15864 4378 15920 4380
rect 15944 4378 16000 4380
rect 16024 4378 16080 4380
rect 16104 4378 16160 4380
rect 15864 4326 15910 4378
rect 15910 4326 15920 4378
rect 15944 4326 15974 4378
rect 15974 4326 15986 4378
rect 15986 4326 16000 4378
rect 16024 4326 16038 4378
rect 16038 4326 16050 4378
rect 16050 4326 16080 4378
rect 16104 4326 16114 4378
rect 16114 4326 16160 4378
rect 15864 4324 15920 4326
rect 15944 4324 16000 4326
rect 16024 4324 16080 4326
rect 16104 4324 16160 4326
rect 15204 3834 15260 3836
rect 15284 3834 15340 3836
rect 15364 3834 15420 3836
rect 15444 3834 15500 3836
rect 15204 3782 15250 3834
rect 15250 3782 15260 3834
rect 15284 3782 15314 3834
rect 15314 3782 15326 3834
rect 15326 3782 15340 3834
rect 15364 3782 15378 3834
rect 15378 3782 15390 3834
rect 15390 3782 15420 3834
rect 15444 3782 15454 3834
rect 15454 3782 15500 3834
rect 15204 3780 15260 3782
rect 15284 3780 15340 3782
rect 15364 3780 15420 3782
rect 15444 3780 15500 3782
rect 17038 10240 17094 10296
rect 17038 8880 17094 8936
rect 17038 7520 17094 7576
rect 17038 6840 17094 6896
rect 15864 3290 15920 3292
rect 15944 3290 16000 3292
rect 16024 3290 16080 3292
rect 16104 3290 16160 3292
rect 15864 3238 15910 3290
rect 15910 3238 15920 3290
rect 15944 3238 15974 3290
rect 15974 3238 15986 3290
rect 15986 3238 16000 3290
rect 16024 3238 16038 3290
rect 16038 3238 16050 3290
rect 16050 3238 16080 3290
rect 16104 3238 16114 3290
rect 16114 3238 16160 3290
rect 15864 3236 15920 3238
rect 15944 3236 16000 3238
rect 16024 3236 16080 3238
rect 16104 3236 16160 3238
rect 17038 5480 17094 5536
rect 17038 3476 17040 3496
rect 17040 3476 17092 3496
rect 17092 3476 17094 3496
rect 17038 3440 17094 3476
rect 17038 2760 17094 2816
rect 15204 2746 15260 2748
rect 15284 2746 15340 2748
rect 15364 2746 15420 2748
rect 15444 2746 15500 2748
rect 15204 2694 15250 2746
rect 15250 2694 15260 2746
rect 15284 2694 15314 2746
rect 15314 2694 15326 2746
rect 15326 2694 15340 2746
rect 15364 2694 15378 2746
rect 15378 2694 15390 2746
rect 15390 2694 15420 2746
rect 15444 2694 15454 2746
rect 15454 2694 15500 2746
rect 15204 2692 15260 2694
rect 15284 2692 15340 2694
rect 15364 2692 15420 2694
rect 15444 2692 15500 2694
rect 3651 2202 3707 2204
rect 3731 2202 3787 2204
rect 3811 2202 3867 2204
rect 3891 2202 3947 2204
rect 3651 2150 3697 2202
rect 3697 2150 3707 2202
rect 3731 2150 3761 2202
rect 3761 2150 3773 2202
rect 3773 2150 3787 2202
rect 3811 2150 3825 2202
rect 3825 2150 3837 2202
rect 3837 2150 3867 2202
rect 3891 2150 3901 2202
rect 3901 2150 3947 2202
rect 3651 2148 3707 2150
rect 3731 2148 3787 2150
rect 3811 2148 3867 2150
rect 3891 2148 3947 2150
rect 7722 2202 7778 2204
rect 7802 2202 7858 2204
rect 7882 2202 7938 2204
rect 7962 2202 8018 2204
rect 7722 2150 7768 2202
rect 7768 2150 7778 2202
rect 7802 2150 7832 2202
rect 7832 2150 7844 2202
rect 7844 2150 7858 2202
rect 7882 2150 7896 2202
rect 7896 2150 7908 2202
rect 7908 2150 7938 2202
rect 7962 2150 7972 2202
rect 7972 2150 8018 2202
rect 7722 2148 7778 2150
rect 7802 2148 7858 2150
rect 7882 2148 7938 2150
rect 7962 2148 8018 2150
rect 11793 2202 11849 2204
rect 11873 2202 11929 2204
rect 11953 2202 12009 2204
rect 12033 2202 12089 2204
rect 11793 2150 11839 2202
rect 11839 2150 11849 2202
rect 11873 2150 11903 2202
rect 11903 2150 11915 2202
rect 11915 2150 11929 2202
rect 11953 2150 11967 2202
rect 11967 2150 11979 2202
rect 11979 2150 12009 2202
rect 12033 2150 12043 2202
rect 12043 2150 12089 2202
rect 11793 2148 11849 2150
rect 11873 2148 11929 2150
rect 11953 2148 12009 2150
rect 12033 2148 12089 2150
rect 15864 2202 15920 2204
rect 15944 2202 16000 2204
rect 16024 2202 16080 2204
rect 16104 2202 16160 2204
rect 15864 2150 15910 2202
rect 15910 2150 15920 2202
rect 15944 2150 15974 2202
rect 15974 2150 15986 2202
rect 15986 2150 16000 2202
rect 16024 2150 16038 2202
rect 16038 2150 16050 2202
rect 16050 2150 16080 2202
rect 16104 2150 16114 2202
rect 16114 2150 16160 2202
rect 15864 2148 15920 2150
rect 15944 2148 16000 2150
rect 16024 2148 16080 2150
rect 16104 2148 16160 2150
<< metal3 >>
rect 2981 17984 3297 17985
rect 2981 17920 2987 17984
rect 3051 17920 3067 17984
rect 3131 17920 3147 17984
rect 3211 17920 3227 17984
rect 3291 17920 3297 17984
rect 2981 17919 3297 17920
rect 7052 17984 7368 17985
rect 7052 17920 7058 17984
rect 7122 17920 7138 17984
rect 7202 17920 7218 17984
rect 7282 17920 7298 17984
rect 7362 17920 7368 17984
rect 7052 17919 7368 17920
rect 11123 17984 11439 17985
rect 11123 17920 11129 17984
rect 11193 17920 11209 17984
rect 11273 17920 11289 17984
rect 11353 17920 11369 17984
rect 11433 17920 11439 17984
rect 11123 17919 11439 17920
rect 15194 17984 15510 17985
rect 15194 17920 15200 17984
rect 15264 17920 15280 17984
rect 15344 17920 15360 17984
rect 15424 17920 15440 17984
rect 15504 17920 15510 17984
rect 15194 17919 15510 17920
rect 3641 17440 3957 17441
rect 3641 17376 3647 17440
rect 3711 17376 3727 17440
rect 3791 17376 3807 17440
rect 3871 17376 3887 17440
rect 3951 17376 3957 17440
rect 3641 17375 3957 17376
rect 7712 17440 8028 17441
rect 7712 17376 7718 17440
rect 7782 17376 7798 17440
rect 7862 17376 7878 17440
rect 7942 17376 7958 17440
rect 8022 17376 8028 17440
rect 7712 17375 8028 17376
rect 11783 17440 12099 17441
rect 11783 17376 11789 17440
rect 11853 17376 11869 17440
rect 11933 17376 11949 17440
rect 12013 17376 12029 17440
rect 12093 17376 12099 17440
rect 11783 17375 12099 17376
rect 15854 17440 16170 17441
rect 15854 17376 15860 17440
rect 15924 17376 15940 17440
rect 16004 17376 16020 17440
rect 16084 17376 16100 17440
rect 16164 17376 16170 17440
rect 15854 17375 16170 17376
rect 841 17234 907 17237
rect 798 17232 907 17234
rect 798 17176 846 17232
rect 902 17176 907 17232
rect 798 17171 907 17176
rect 798 17128 858 17171
rect 0 17038 858 17128
rect 0 17008 800 17038
rect 2981 16896 3297 16897
rect 2981 16832 2987 16896
rect 3051 16832 3067 16896
rect 3131 16832 3147 16896
rect 3211 16832 3227 16896
rect 3291 16832 3297 16896
rect 2981 16831 3297 16832
rect 7052 16896 7368 16897
rect 7052 16832 7058 16896
rect 7122 16832 7138 16896
rect 7202 16832 7218 16896
rect 7282 16832 7298 16896
rect 7362 16832 7368 16896
rect 7052 16831 7368 16832
rect 11123 16896 11439 16897
rect 11123 16832 11129 16896
rect 11193 16832 11209 16896
rect 11273 16832 11289 16896
rect 11353 16832 11369 16896
rect 11433 16832 11439 16896
rect 11123 16831 11439 16832
rect 15194 16896 15510 16897
rect 15194 16832 15200 16896
rect 15264 16832 15280 16896
rect 15344 16832 15360 16896
rect 15424 16832 15440 16896
rect 15504 16832 15510 16896
rect 15194 16831 15510 16832
rect 3641 16352 3957 16353
rect 3641 16288 3647 16352
rect 3711 16288 3727 16352
rect 3791 16288 3807 16352
rect 3871 16288 3887 16352
rect 3951 16288 3957 16352
rect 3641 16287 3957 16288
rect 7712 16352 8028 16353
rect 7712 16288 7718 16352
rect 7782 16288 7798 16352
rect 7862 16288 7878 16352
rect 7942 16288 7958 16352
rect 8022 16288 8028 16352
rect 7712 16287 8028 16288
rect 11783 16352 12099 16353
rect 11783 16288 11789 16352
rect 11853 16288 11869 16352
rect 11933 16288 11949 16352
rect 12013 16288 12029 16352
rect 12093 16288 12099 16352
rect 11783 16287 12099 16288
rect 15854 16352 16170 16353
rect 15854 16288 15860 16352
rect 15924 16288 15940 16352
rect 16004 16288 16020 16352
rect 16084 16288 16100 16352
rect 16164 16288 16170 16352
rect 15854 16287 16170 16288
rect 2981 15808 3297 15809
rect 0 15738 800 15768
rect 2981 15744 2987 15808
rect 3051 15744 3067 15808
rect 3131 15744 3147 15808
rect 3211 15744 3227 15808
rect 3291 15744 3297 15808
rect 2981 15743 3297 15744
rect 7052 15808 7368 15809
rect 7052 15744 7058 15808
rect 7122 15744 7138 15808
rect 7202 15744 7218 15808
rect 7282 15744 7298 15808
rect 7362 15744 7368 15808
rect 7052 15743 7368 15744
rect 11123 15808 11439 15809
rect 11123 15744 11129 15808
rect 11193 15744 11209 15808
rect 11273 15744 11289 15808
rect 11353 15744 11369 15808
rect 11433 15744 11439 15808
rect 11123 15743 11439 15744
rect 15194 15808 15510 15809
rect 15194 15744 15200 15808
rect 15264 15744 15280 15808
rect 15344 15744 15360 15808
rect 15424 15744 15440 15808
rect 15504 15744 15510 15808
rect 15194 15743 15510 15744
rect 1025 15738 1091 15741
rect 0 15736 1091 15738
rect 0 15680 1030 15736
rect 1086 15680 1091 15736
rect 0 15678 1091 15680
rect 0 15648 800 15678
rect 1025 15675 1091 15678
rect 3641 15264 3957 15265
rect 3641 15200 3647 15264
rect 3711 15200 3727 15264
rect 3791 15200 3807 15264
rect 3871 15200 3887 15264
rect 3951 15200 3957 15264
rect 3641 15199 3957 15200
rect 7712 15264 8028 15265
rect 7712 15200 7718 15264
rect 7782 15200 7798 15264
rect 7862 15200 7878 15264
rect 7942 15200 7958 15264
rect 8022 15200 8028 15264
rect 7712 15199 8028 15200
rect 11783 15264 12099 15265
rect 11783 15200 11789 15264
rect 11853 15200 11869 15264
rect 11933 15200 11949 15264
rect 12013 15200 12029 15264
rect 12093 15200 12099 15264
rect 11783 15199 12099 15200
rect 15854 15264 16170 15265
rect 15854 15200 15860 15264
rect 15924 15200 15940 15264
rect 16004 15200 16020 15264
rect 16084 15200 16100 15264
rect 16164 15200 16170 15264
rect 15854 15199 16170 15200
rect 16849 15058 16915 15061
rect 17716 15058 18516 15088
rect 16849 15056 18516 15058
rect 16849 15000 16854 15056
rect 16910 15000 18516 15056
rect 16849 14998 18516 15000
rect 16849 14995 16915 14998
rect 17716 14968 18516 14998
rect 2981 14720 3297 14721
rect 2981 14656 2987 14720
rect 3051 14656 3067 14720
rect 3131 14656 3147 14720
rect 3211 14656 3227 14720
rect 3291 14656 3297 14720
rect 2981 14655 3297 14656
rect 7052 14720 7368 14721
rect 7052 14656 7058 14720
rect 7122 14656 7138 14720
rect 7202 14656 7218 14720
rect 7282 14656 7298 14720
rect 7362 14656 7368 14720
rect 7052 14655 7368 14656
rect 11123 14720 11439 14721
rect 11123 14656 11129 14720
rect 11193 14656 11209 14720
rect 11273 14656 11289 14720
rect 11353 14656 11369 14720
rect 11433 14656 11439 14720
rect 11123 14655 11439 14656
rect 15194 14720 15510 14721
rect 15194 14656 15200 14720
rect 15264 14656 15280 14720
rect 15344 14656 15360 14720
rect 15424 14656 15440 14720
rect 15504 14656 15510 14720
rect 15194 14655 15510 14656
rect 17033 14378 17099 14381
rect 17716 14378 18516 14408
rect 17033 14376 18516 14378
rect 17033 14320 17038 14376
rect 17094 14320 18516 14376
rect 17033 14318 18516 14320
rect 17033 14315 17099 14318
rect 17716 14288 18516 14318
rect 3641 14176 3957 14177
rect 3641 14112 3647 14176
rect 3711 14112 3727 14176
rect 3791 14112 3807 14176
rect 3871 14112 3887 14176
rect 3951 14112 3957 14176
rect 3641 14111 3957 14112
rect 7712 14176 8028 14177
rect 7712 14112 7718 14176
rect 7782 14112 7798 14176
rect 7862 14112 7878 14176
rect 7942 14112 7958 14176
rect 8022 14112 8028 14176
rect 7712 14111 8028 14112
rect 11783 14176 12099 14177
rect 11783 14112 11789 14176
rect 11853 14112 11869 14176
rect 11933 14112 11949 14176
rect 12013 14112 12029 14176
rect 12093 14112 12099 14176
rect 11783 14111 12099 14112
rect 15854 14176 16170 14177
rect 15854 14112 15860 14176
rect 15924 14112 15940 14176
rect 16004 14112 16020 14176
rect 16084 14112 16100 14176
rect 16164 14112 16170 14176
rect 15854 14111 16170 14112
rect 0 13698 800 13728
rect 1393 13698 1459 13701
rect 0 13696 1459 13698
rect 0 13640 1398 13696
rect 1454 13640 1459 13696
rect 0 13638 1459 13640
rect 0 13608 800 13638
rect 1393 13635 1459 13638
rect 2981 13632 3297 13633
rect 2981 13568 2987 13632
rect 3051 13568 3067 13632
rect 3131 13568 3147 13632
rect 3211 13568 3227 13632
rect 3291 13568 3297 13632
rect 2981 13567 3297 13568
rect 7052 13632 7368 13633
rect 7052 13568 7058 13632
rect 7122 13568 7138 13632
rect 7202 13568 7218 13632
rect 7282 13568 7298 13632
rect 7362 13568 7368 13632
rect 7052 13567 7368 13568
rect 11123 13632 11439 13633
rect 11123 13568 11129 13632
rect 11193 13568 11209 13632
rect 11273 13568 11289 13632
rect 11353 13568 11369 13632
rect 11433 13568 11439 13632
rect 11123 13567 11439 13568
rect 15194 13632 15510 13633
rect 15194 13568 15200 13632
rect 15264 13568 15280 13632
rect 15344 13568 15360 13632
rect 15424 13568 15440 13632
rect 15504 13568 15510 13632
rect 15194 13567 15510 13568
rect 841 13154 907 13157
rect 798 13152 907 13154
rect 798 13096 846 13152
rect 902 13096 907 13152
rect 798 13091 907 13096
rect 798 13048 858 13091
rect 0 12958 858 13048
rect 3641 13088 3957 13089
rect 3641 13024 3647 13088
rect 3711 13024 3727 13088
rect 3791 13024 3807 13088
rect 3871 13024 3887 13088
rect 3951 13024 3957 13088
rect 3641 13023 3957 13024
rect 7712 13088 8028 13089
rect 7712 13024 7718 13088
rect 7782 13024 7798 13088
rect 7862 13024 7878 13088
rect 7942 13024 7958 13088
rect 8022 13024 8028 13088
rect 7712 13023 8028 13024
rect 11783 13088 12099 13089
rect 11783 13024 11789 13088
rect 11853 13024 11869 13088
rect 11933 13024 11949 13088
rect 12013 13024 12029 13088
rect 12093 13024 12099 13088
rect 11783 13023 12099 13024
rect 15854 13088 16170 13089
rect 15854 13024 15860 13088
rect 15924 13024 15940 13088
rect 16004 13024 16020 13088
rect 16084 13024 16100 13088
rect 16164 13024 16170 13088
rect 15854 13023 16170 13024
rect 17033 13018 17099 13021
rect 17716 13018 18516 13048
rect 17033 13016 18516 13018
rect 17033 12960 17038 13016
rect 17094 12960 18516 13016
rect 17033 12958 18516 12960
rect 0 12928 800 12958
rect 17033 12955 17099 12958
rect 17716 12928 18516 12958
rect 2981 12544 3297 12545
rect 2981 12480 2987 12544
rect 3051 12480 3067 12544
rect 3131 12480 3147 12544
rect 3211 12480 3227 12544
rect 3291 12480 3297 12544
rect 2981 12479 3297 12480
rect 7052 12544 7368 12545
rect 7052 12480 7058 12544
rect 7122 12480 7138 12544
rect 7202 12480 7218 12544
rect 7282 12480 7298 12544
rect 7362 12480 7368 12544
rect 7052 12479 7368 12480
rect 11123 12544 11439 12545
rect 11123 12480 11129 12544
rect 11193 12480 11209 12544
rect 11273 12480 11289 12544
rect 11353 12480 11369 12544
rect 11433 12480 11439 12544
rect 11123 12479 11439 12480
rect 15194 12544 15510 12545
rect 15194 12480 15200 12544
rect 15264 12480 15280 12544
rect 15344 12480 15360 12544
rect 15424 12480 15440 12544
rect 15504 12480 15510 12544
rect 15194 12479 15510 12480
rect 3641 12000 3957 12001
rect 3641 11936 3647 12000
rect 3711 11936 3727 12000
rect 3791 11936 3807 12000
rect 3871 11936 3887 12000
rect 3951 11936 3957 12000
rect 3641 11935 3957 11936
rect 7712 12000 8028 12001
rect 7712 11936 7718 12000
rect 7782 11936 7798 12000
rect 7862 11936 7878 12000
rect 7942 11936 7958 12000
rect 8022 11936 8028 12000
rect 7712 11935 8028 11936
rect 11783 12000 12099 12001
rect 11783 11936 11789 12000
rect 11853 11936 11869 12000
rect 11933 11936 11949 12000
rect 12013 11936 12029 12000
rect 12093 11936 12099 12000
rect 11783 11935 12099 11936
rect 15854 12000 16170 12001
rect 15854 11936 15860 12000
rect 15924 11936 15940 12000
rect 16004 11936 16020 12000
rect 16084 11936 16100 12000
rect 16164 11936 16170 12000
rect 15854 11935 16170 11936
rect 16481 11658 16547 11661
rect 17716 11658 18516 11688
rect 16481 11656 18516 11658
rect 16481 11600 16486 11656
rect 16542 11600 18516 11656
rect 16481 11598 18516 11600
rect 16481 11595 16547 11598
rect 17716 11568 18516 11598
rect 2981 11456 3297 11457
rect 2981 11392 2987 11456
rect 3051 11392 3067 11456
rect 3131 11392 3147 11456
rect 3211 11392 3227 11456
rect 3291 11392 3297 11456
rect 2981 11391 3297 11392
rect 7052 11456 7368 11457
rect 7052 11392 7058 11456
rect 7122 11392 7138 11456
rect 7202 11392 7218 11456
rect 7282 11392 7298 11456
rect 7362 11392 7368 11456
rect 7052 11391 7368 11392
rect 11123 11456 11439 11457
rect 11123 11392 11129 11456
rect 11193 11392 11209 11456
rect 11273 11392 11289 11456
rect 11353 11392 11369 11456
rect 11433 11392 11439 11456
rect 11123 11391 11439 11392
rect 15194 11456 15510 11457
rect 15194 11392 15200 11456
rect 15264 11392 15280 11456
rect 15344 11392 15360 11456
rect 15424 11392 15440 11456
rect 15504 11392 15510 11456
rect 15194 11391 15510 11392
rect 0 10978 800 11008
rect 17033 10978 17099 10981
rect 17716 10978 18516 11008
rect 0 10888 858 10978
rect 17033 10976 18516 10978
rect 17033 10920 17038 10976
rect 17094 10920 18516 10976
rect 17033 10918 18516 10920
rect 17033 10915 17099 10918
rect 798 10845 858 10888
rect 3641 10912 3957 10913
rect 3641 10848 3647 10912
rect 3711 10848 3727 10912
rect 3791 10848 3807 10912
rect 3871 10848 3887 10912
rect 3951 10848 3957 10912
rect 3641 10847 3957 10848
rect 7712 10912 8028 10913
rect 7712 10848 7718 10912
rect 7782 10848 7798 10912
rect 7862 10848 7878 10912
rect 7942 10848 7958 10912
rect 8022 10848 8028 10912
rect 7712 10847 8028 10848
rect 11783 10912 12099 10913
rect 11783 10848 11789 10912
rect 11853 10848 11869 10912
rect 11933 10848 11949 10912
rect 12013 10848 12029 10912
rect 12093 10848 12099 10912
rect 11783 10847 12099 10848
rect 15854 10912 16170 10913
rect 15854 10848 15860 10912
rect 15924 10848 15940 10912
rect 16004 10848 16020 10912
rect 16084 10848 16100 10912
rect 16164 10848 16170 10912
rect 17716 10888 18516 10918
rect 15854 10847 16170 10848
rect 798 10840 907 10845
rect 798 10784 846 10840
rect 902 10784 907 10840
rect 798 10782 907 10784
rect 841 10779 907 10782
rect 2981 10368 3297 10369
rect 2981 10304 2987 10368
rect 3051 10304 3067 10368
rect 3131 10304 3147 10368
rect 3211 10304 3227 10368
rect 3291 10304 3297 10368
rect 2981 10303 3297 10304
rect 7052 10368 7368 10369
rect 7052 10304 7058 10368
rect 7122 10304 7138 10368
rect 7202 10304 7218 10368
rect 7282 10304 7298 10368
rect 7362 10304 7368 10368
rect 7052 10303 7368 10304
rect 11123 10368 11439 10369
rect 11123 10304 11129 10368
rect 11193 10304 11209 10368
rect 11273 10304 11289 10368
rect 11353 10304 11369 10368
rect 11433 10304 11439 10368
rect 11123 10303 11439 10304
rect 15194 10368 15510 10369
rect 15194 10304 15200 10368
rect 15264 10304 15280 10368
rect 15344 10304 15360 10368
rect 15424 10304 15440 10368
rect 15504 10304 15510 10368
rect 15194 10303 15510 10304
rect 17033 10298 17099 10301
rect 17716 10298 18516 10328
rect 17033 10296 18516 10298
rect 17033 10240 17038 10296
rect 17094 10240 18516 10296
rect 17033 10238 18516 10240
rect 17033 10235 17099 10238
rect 17716 10208 18516 10238
rect 3641 9824 3957 9825
rect 3641 9760 3647 9824
rect 3711 9760 3727 9824
rect 3791 9760 3807 9824
rect 3871 9760 3887 9824
rect 3951 9760 3957 9824
rect 3641 9759 3957 9760
rect 7712 9824 8028 9825
rect 7712 9760 7718 9824
rect 7782 9760 7798 9824
rect 7862 9760 7878 9824
rect 7942 9760 7958 9824
rect 8022 9760 8028 9824
rect 7712 9759 8028 9760
rect 11783 9824 12099 9825
rect 11783 9760 11789 9824
rect 11853 9760 11869 9824
rect 11933 9760 11949 9824
rect 12013 9760 12029 9824
rect 12093 9760 12099 9824
rect 11783 9759 12099 9760
rect 15854 9824 16170 9825
rect 15854 9760 15860 9824
rect 15924 9760 15940 9824
rect 16004 9760 16020 9824
rect 16084 9760 16100 9824
rect 16164 9760 16170 9824
rect 15854 9759 16170 9760
rect 0 9618 800 9648
rect 1393 9618 1459 9621
rect 0 9616 1459 9618
rect 0 9560 1398 9616
rect 1454 9560 1459 9616
rect 0 9558 1459 9560
rect 0 9528 800 9558
rect 1393 9555 1459 9558
rect 2957 9618 3023 9621
rect 3417 9618 3483 9621
rect 2957 9616 3483 9618
rect 2957 9560 2962 9616
rect 3018 9560 3422 9616
rect 3478 9560 3483 9616
rect 2957 9558 3483 9560
rect 2957 9555 3023 9558
rect 3417 9555 3483 9558
rect 2405 9482 2471 9485
rect 3325 9482 3391 9485
rect 2405 9480 3391 9482
rect 2405 9424 2410 9480
rect 2466 9424 3330 9480
rect 3386 9424 3391 9480
rect 2405 9422 3391 9424
rect 2405 9419 2471 9422
rect 3325 9419 3391 9422
rect 2981 9280 3297 9281
rect 2981 9216 2987 9280
rect 3051 9216 3067 9280
rect 3131 9216 3147 9280
rect 3211 9216 3227 9280
rect 3291 9216 3297 9280
rect 2981 9215 3297 9216
rect 7052 9280 7368 9281
rect 7052 9216 7058 9280
rect 7122 9216 7138 9280
rect 7202 9216 7218 9280
rect 7282 9216 7298 9280
rect 7362 9216 7368 9280
rect 7052 9215 7368 9216
rect 11123 9280 11439 9281
rect 11123 9216 11129 9280
rect 11193 9216 11209 9280
rect 11273 9216 11289 9280
rect 11353 9216 11369 9280
rect 11433 9216 11439 9280
rect 11123 9215 11439 9216
rect 15194 9280 15510 9281
rect 15194 9216 15200 9280
rect 15264 9216 15280 9280
rect 15344 9216 15360 9280
rect 15424 9216 15440 9280
rect 15504 9216 15510 9280
rect 15194 9215 15510 9216
rect 0 8938 800 8968
rect 17033 8938 17099 8941
rect 17716 8938 18516 8968
rect 0 8848 858 8938
rect 17033 8936 18516 8938
rect 17033 8880 17038 8936
rect 17094 8880 18516 8936
rect 17033 8878 18516 8880
rect 17033 8875 17099 8878
rect 17716 8848 18516 8878
rect 798 8805 858 8848
rect 798 8800 907 8805
rect 798 8744 846 8800
rect 902 8744 907 8800
rect 798 8742 907 8744
rect 841 8739 907 8742
rect 3641 8736 3957 8737
rect 3641 8672 3647 8736
rect 3711 8672 3727 8736
rect 3791 8672 3807 8736
rect 3871 8672 3887 8736
rect 3951 8672 3957 8736
rect 3641 8671 3957 8672
rect 7712 8736 8028 8737
rect 7712 8672 7718 8736
rect 7782 8672 7798 8736
rect 7862 8672 7878 8736
rect 7942 8672 7958 8736
rect 8022 8672 8028 8736
rect 7712 8671 8028 8672
rect 11783 8736 12099 8737
rect 11783 8672 11789 8736
rect 11853 8672 11869 8736
rect 11933 8672 11949 8736
rect 12013 8672 12029 8736
rect 12093 8672 12099 8736
rect 11783 8671 12099 8672
rect 15854 8736 16170 8737
rect 15854 8672 15860 8736
rect 15924 8672 15940 8736
rect 16004 8672 16020 8736
rect 16084 8672 16100 8736
rect 16164 8672 16170 8736
rect 15854 8671 16170 8672
rect 0 8258 800 8288
rect 1669 8258 1735 8261
rect 0 8256 1735 8258
rect 0 8200 1674 8256
rect 1730 8200 1735 8256
rect 0 8198 1735 8200
rect 0 8168 800 8198
rect 1669 8195 1735 8198
rect 2981 8192 3297 8193
rect 2981 8128 2987 8192
rect 3051 8128 3067 8192
rect 3131 8128 3147 8192
rect 3211 8128 3227 8192
rect 3291 8128 3297 8192
rect 2981 8127 3297 8128
rect 7052 8192 7368 8193
rect 7052 8128 7058 8192
rect 7122 8128 7138 8192
rect 7202 8128 7218 8192
rect 7282 8128 7298 8192
rect 7362 8128 7368 8192
rect 7052 8127 7368 8128
rect 11123 8192 11439 8193
rect 11123 8128 11129 8192
rect 11193 8128 11209 8192
rect 11273 8128 11289 8192
rect 11353 8128 11369 8192
rect 11433 8128 11439 8192
rect 11123 8127 11439 8128
rect 15194 8192 15510 8193
rect 15194 8128 15200 8192
rect 15264 8128 15280 8192
rect 15344 8128 15360 8192
rect 15424 8128 15440 8192
rect 15504 8128 15510 8192
rect 15194 8127 15510 8128
rect 841 7714 907 7717
rect 798 7712 907 7714
rect 798 7656 846 7712
rect 902 7656 907 7712
rect 798 7651 907 7656
rect 798 7608 858 7651
rect 0 7518 858 7608
rect 3641 7648 3957 7649
rect 3641 7584 3647 7648
rect 3711 7584 3727 7648
rect 3791 7584 3807 7648
rect 3871 7584 3887 7648
rect 3951 7584 3957 7648
rect 3641 7583 3957 7584
rect 7712 7648 8028 7649
rect 7712 7584 7718 7648
rect 7782 7584 7798 7648
rect 7862 7584 7878 7648
rect 7942 7584 7958 7648
rect 8022 7584 8028 7648
rect 7712 7583 8028 7584
rect 11783 7648 12099 7649
rect 11783 7584 11789 7648
rect 11853 7584 11869 7648
rect 11933 7584 11949 7648
rect 12013 7584 12029 7648
rect 12093 7584 12099 7648
rect 11783 7583 12099 7584
rect 15854 7648 16170 7649
rect 15854 7584 15860 7648
rect 15924 7584 15940 7648
rect 16004 7584 16020 7648
rect 16084 7584 16100 7648
rect 16164 7584 16170 7648
rect 15854 7583 16170 7584
rect 17033 7578 17099 7581
rect 17716 7578 18516 7608
rect 17033 7576 18516 7578
rect 17033 7520 17038 7576
rect 17094 7520 18516 7576
rect 17033 7518 18516 7520
rect 0 7488 800 7518
rect 17033 7515 17099 7518
rect 17716 7488 18516 7518
rect 2981 7104 3297 7105
rect 2981 7040 2987 7104
rect 3051 7040 3067 7104
rect 3131 7040 3147 7104
rect 3211 7040 3227 7104
rect 3291 7040 3297 7104
rect 2981 7039 3297 7040
rect 7052 7104 7368 7105
rect 7052 7040 7058 7104
rect 7122 7040 7138 7104
rect 7202 7040 7218 7104
rect 7282 7040 7298 7104
rect 7362 7040 7368 7104
rect 7052 7039 7368 7040
rect 11123 7104 11439 7105
rect 11123 7040 11129 7104
rect 11193 7040 11209 7104
rect 11273 7040 11289 7104
rect 11353 7040 11369 7104
rect 11433 7040 11439 7104
rect 11123 7039 11439 7040
rect 15194 7104 15510 7105
rect 15194 7040 15200 7104
rect 15264 7040 15280 7104
rect 15344 7040 15360 7104
rect 15424 7040 15440 7104
rect 15504 7040 15510 7104
rect 15194 7039 15510 7040
rect 0 6898 800 6928
rect 4061 6898 4127 6901
rect 0 6896 4127 6898
rect 0 6840 4066 6896
rect 4122 6840 4127 6896
rect 0 6838 4127 6840
rect 0 6808 800 6838
rect 4061 6835 4127 6838
rect 17033 6898 17099 6901
rect 17716 6898 18516 6928
rect 17033 6896 18516 6898
rect 17033 6840 17038 6896
rect 17094 6840 18516 6896
rect 17033 6838 18516 6840
rect 17033 6835 17099 6838
rect 17716 6808 18516 6838
rect 3641 6560 3957 6561
rect 3641 6496 3647 6560
rect 3711 6496 3727 6560
rect 3791 6496 3807 6560
rect 3871 6496 3887 6560
rect 3951 6496 3957 6560
rect 3641 6495 3957 6496
rect 7712 6560 8028 6561
rect 7712 6496 7718 6560
rect 7782 6496 7798 6560
rect 7862 6496 7878 6560
rect 7942 6496 7958 6560
rect 8022 6496 8028 6560
rect 7712 6495 8028 6496
rect 11783 6560 12099 6561
rect 11783 6496 11789 6560
rect 11853 6496 11869 6560
rect 11933 6496 11949 6560
rect 12013 6496 12029 6560
rect 12093 6496 12099 6560
rect 11783 6495 12099 6496
rect 15854 6560 16170 6561
rect 15854 6496 15860 6560
rect 15924 6496 15940 6560
rect 16004 6496 16020 6560
rect 16084 6496 16100 6560
rect 16164 6496 16170 6560
rect 15854 6495 16170 6496
rect 2981 6016 3297 6017
rect 2981 5952 2987 6016
rect 3051 5952 3067 6016
rect 3131 5952 3147 6016
rect 3211 5952 3227 6016
rect 3291 5952 3297 6016
rect 2981 5951 3297 5952
rect 7052 6016 7368 6017
rect 7052 5952 7058 6016
rect 7122 5952 7138 6016
rect 7202 5952 7218 6016
rect 7282 5952 7298 6016
rect 7362 5952 7368 6016
rect 7052 5951 7368 5952
rect 11123 6016 11439 6017
rect 11123 5952 11129 6016
rect 11193 5952 11209 6016
rect 11273 5952 11289 6016
rect 11353 5952 11369 6016
rect 11433 5952 11439 6016
rect 11123 5951 11439 5952
rect 15194 6016 15510 6017
rect 15194 5952 15200 6016
rect 15264 5952 15280 6016
rect 15344 5952 15360 6016
rect 15424 5952 15440 6016
rect 15504 5952 15510 6016
rect 15194 5951 15510 5952
rect 0 5538 800 5568
rect 1393 5538 1459 5541
rect 0 5536 1459 5538
rect 0 5480 1398 5536
rect 1454 5480 1459 5536
rect 0 5478 1459 5480
rect 0 5448 800 5478
rect 1393 5475 1459 5478
rect 17033 5538 17099 5541
rect 17716 5538 18516 5568
rect 17033 5536 18516 5538
rect 17033 5480 17038 5536
rect 17094 5480 18516 5536
rect 17033 5478 18516 5480
rect 17033 5475 17099 5478
rect 3641 5472 3957 5473
rect 3641 5408 3647 5472
rect 3711 5408 3727 5472
rect 3791 5408 3807 5472
rect 3871 5408 3887 5472
rect 3951 5408 3957 5472
rect 3641 5407 3957 5408
rect 7712 5472 8028 5473
rect 7712 5408 7718 5472
rect 7782 5408 7798 5472
rect 7862 5408 7878 5472
rect 7942 5408 7958 5472
rect 8022 5408 8028 5472
rect 7712 5407 8028 5408
rect 11783 5472 12099 5473
rect 11783 5408 11789 5472
rect 11853 5408 11869 5472
rect 11933 5408 11949 5472
rect 12013 5408 12029 5472
rect 12093 5408 12099 5472
rect 11783 5407 12099 5408
rect 15854 5472 16170 5473
rect 15854 5408 15860 5472
rect 15924 5408 15940 5472
rect 16004 5408 16020 5472
rect 16084 5408 16100 5472
rect 16164 5408 16170 5472
rect 17716 5448 18516 5478
rect 15854 5407 16170 5408
rect 2981 4928 3297 4929
rect 2981 4864 2987 4928
rect 3051 4864 3067 4928
rect 3131 4864 3147 4928
rect 3211 4864 3227 4928
rect 3291 4864 3297 4928
rect 2981 4863 3297 4864
rect 7052 4928 7368 4929
rect 7052 4864 7058 4928
rect 7122 4864 7138 4928
rect 7202 4864 7218 4928
rect 7282 4864 7298 4928
rect 7362 4864 7368 4928
rect 7052 4863 7368 4864
rect 11123 4928 11439 4929
rect 11123 4864 11129 4928
rect 11193 4864 11209 4928
rect 11273 4864 11289 4928
rect 11353 4864 11369 4928
rect 11433 4864 11439 4928
rect 11123 4863 11439 4864
rect 15194 4928 15510 4929
rect 15194 4864 15200 4928
rect 15264 4864 15280 4928
rect 15344 4864 15360 4928
rect 15424 4864 15440 4928
rect 15504 4864 15510 4928
rect 15194 4863 15510 4864
rect 3641 4384 3957 4385
rect 3641 4320 3647 4384
rect 3711 4320 3727 4384
rect 3791 4320 3807 4384
rect 3871 4320 3887 4384
rect 3951 4320 3957 4384
rect 3641 4319 3957 4320
rect 7712 4384 8028 4385
rect 7712 4320 7718 4384
rect 7782 4320 7798 4384
rect 7862 4320 7878 4384
rect 7942 4320 7958 4384
rect 8022 4320 8028 4384
rect 7712 4319 8028 4320
rect 11783 4384 12099 4385
rect 11783 4320 11789 4384
rect 11853 4320 11869 4384
rect 11933 4320 11949 4384
rect 12013 4320 12029 4384
rect 12093 4320 12099 4384
rect 11783 4319 12099 4320
rect 15854 4384 16170 4385
rect 15854 4320 15860 4384
rect 15924 4320 15940 4384
rect 16004 4320 16020 4384
rect 16084 4320 16100 4384
rect 16164 4320 16170 4384
rect 15854 4319 16170 4320
rect 2981 3840 3297 3841
rect 2981 3776 2987 3840
rect 3051 3776 3067 3840
rect 3131 3776 3147 3840
rect 3211 3776 3227 3840
rect 3291 3776 3297 3840
rect 2981 3775 3297 3776
rect 7052 3840 7368 3841
rect 7052 3776 7058 3840
rect 7122 3776 7138 3840
rect 7202 3776 7218 3840
rect 7282 3776 7298 3840
rect 7362 3776 7368 3840
rect 7052 3775 7368 3776
rect 11123 3840 11439 3841
rect 11123 3776 11129 3840
rect 11193 3776 11209 3840
rect 11273 3776 11289 3840
rect 11353 3776 11369 3840
rect 11433 3776 11439 3840
rect 11123 3775 11439 3776
rect 15194 3840 15510 3841
rect 15194 3776 15200 3840
rect 15264 3776 15280 3840
rect 15344 3776 15360 3840
rect 15424 3776 15440 3840
rect 15504 3776 15510 3840
rect 15194 3775 15510 3776
rect 17033 3498 17099 3501
rect 17716 3498 18516 3528
rect 17033 3496 18516 3498
rect 17033 3440 17038 3496
rect 17094 3440 18516 3496
rect 17033 3438 18516 3440
rect 17033 3435 17099 3438
rect 17716 3408 18516 3438
rect 3641 3296 3957 3297
rect 3641 3232 3647 3296
rect 3711 3232 3727 3296
rect 3791 3232 3807 3296
rect 3871 3232 3887 3296
rect 3951 3232 3957 3296
rect 3641 3231 3957 3232
rect 7712 3296 8028 3297
rect 7712 3232 7718 3296
rect 7782 3232 7798 3296
rect 7862 3232 7878 3296
rect 7942 3232 7958 3296
rect 8022 3232 8028 3296
rect 7712 3231 8028 3232
rect 11783 3296 12099 3297
rect 11783 3232 11789 3296
rect 11853 3232 11869 3296
rect 11933 3232 11949 3296
rect 12013 3232 12029 3296
rect 12093 3232 12099 3296
rect 11783 3231 12099 3232
rect 15854 3296 16170 3297
rect 15854 3232 15860 3296
rect 15924 3232 15940 3296
rect 16004 3232 16020 3296
rect 16084 3232 16100 3296
rect 16164 3232 16170 3296
rect 15854 3231 16170 3232
rect 17033 2818 17099 2821
rect 17716 2818 18516 2848
rect 17033 2816 18516 2818
rect 17033 2760 17038 2816
rect 17094 2760 18516 2816
rect 17033 2758 18516 2760
rect 17033 2755 17099 2758
rect 2981 2752 3297 2753
rect 2981 2688 2987 2752
rect 3051 2688 3067 2752
rect 3131 2688 3147 2752
rect 3211 2688 3227 2752
rect 3291 2688 3297 2752
rect 2981 2687 3297 2688
rect 7052 2752 7368 2753
rect 7052 2688 7058 2752
rect 7122 2688 7138 2752
rect 7202 2688 7218 2752
rect 7282 2688 7298 2752
rect 7362 2688 7368 2752
rect 7052 2687 7368 2688
rect 11123 2752 11439 2753
rect 11123 2688 11129 2752
rect 11193 2688 11209 2752
rect 11273 2688 11289 2752
rect 11353 2688 11369 2752
rect 11433 2688 11439 2752
rect 11123 2687 11439 2688
rect 15194 2752 15510 2753
rect 15194 2688 15200 2752
rect 15264 2688 15280 2752
rect 15344 2688 15360 2752
rect 15424 2688 15440 2752
rect 15504 2688 15510 2752
rect 17716 2728 18516 2758
rect 15194 2687 15510 2688
rect 3641 2208 3957 2209
rect 3641 2144 3647 2208
rect 3711 2144 3727 2208
rect 3791 2144 3807 2208
rect 3871 2144 3887 2208
rect 3951 2144 3957 2208
rect 3641 2143 3957 2144
rect 7712 2208 8028 2209
rect 7712 2144 7718 2208
rect 7782 2144 7798 2208
rect 7862 2144 7878 2208
rect 7942 2144 7958 2208
rect 8022 2144 8028 2208
rect 7712 2143 8028 2144
rect 11783 2208 12099 2209
rect 11783 2144 11789 2208
rect 11853 2144 11869 2208
rect 11933 2144 11949 2208
rect 12013 2144 12029 2208
rect 12093 2144 12099 2208
rect 11783 2143 12099 2144
rect 15854 2208 16170 2209
rect 15854 2144 15860 2208
rect 15924 2144 15940 2208
rect 16004 2144 16020 2208
rect 16084 2144 16100 2208
rect 16164 2144 16170 2208
rect 15854 2143 16170 2144
<< via3 >>
rect 2987 17980 3051 17984
rect 2987 17924 2991 17980
rect 2991 17924 3047 17980
rect 3047 17924 3051 17980
rect 2987 17920 3051 17924
rect 3067 17980 3131 17984
rect 3067 17924 3071 17980
rect 3071 17924 3127 17980
rect 3127 17924 3131 17980
rect 3067 17920 3131 17924
rect 3147 17980 3211 17984
rect 3147 17924 3151 17980
rect 3151 17924 3207 17980
rect 3207 17924 3211 17980
rect 3147 17920 3211 17924
rect 3227 17980 3291 17984
rect 3227 17924 3231 17980
rect 3231 17924 3287 17980
rect 3287 17924 3291 17980
rect 3227 17920 3291 17924
rect 7058 17980 7122 17984
rect 7058 17924 7062 17980
rect 7062 17924 7118 17980
rect 7118 17924 7122 17980
rect 7058 17920 7122 17924
rect 7138 17980 7202 17984
rect 7138 17924 7142 17980
rect 7142 17924 7198 17980
rect 7198 17924 7202 17980
rect 7138 17920 7202 17924
rect 7218 17980 7282 17984
rect 7218 17924 7222 17980
rect 7222 17924 7278 17980
rect 7278 17924 7282 17980
rect 7218 17920 7282 17924
rect 7298 17980 7362 17984
rect 7298 17924 7302 17980
rect 7302 17924 7358 17980
rect 7358 17924 7362 17980
rect 7298 17920 7362 17924
rect 11129 17980 11193 17984
rect 11129 17924 11133 17980
rect 11133 17924 11189 17980
rect 11189 17924 11193 17980
rect 11129 17920 11193 17924
rect 11209 17980 11273 17984
rect 11209 17924 11213 17980
rect 11213 17924 11269 17980
rect 11269 17924 11273 17980
rect 11209 17920 11273 17924
rect 11289 17980 11353 17984
rect 11289 17924 11293 17980
rect 11293 17924 11349 17980
rect 11349 17924 11353 17980
rect 11289 17920 11353 17924
rect 11369 17980 11433 17984
rect 11369 17924 11373 17980
rect 11373 17924 11429 17980
rect 11429 17924 11433 17980
rect 11369 17920 11433 17924
rect 15200 17980 15264 17984
rect 15200 17924 15204 17980
rect 15204 17924 15260 17980
rect 15260 17924 15264 17980
rect 15200 17920 15264 17924
rect 15280 17980 15344 17984
rect 15280 17924 15284 17980
rect 15284 17924 15340 17980
rect 15340 17924 15344 17980
rect 15280 17920 15344 17924
rect 15360 17980 15424 17984
rect 15360 17924 15364 17980
rect 15364 17924 15420 17980
rect 15420 17924 15424 17980
rect 15360 17920 15424 17924
rect 15440 17980 15504 17984
rect 15440 17924 15444 17980
rect 15444 17924 15500 17980
rect 15500 17924 15504 17980
rect 15440 17920 15504 17924
rect 3647 17436 3711 17440
rect 3647 17380 3651 17436
rect 3651 17380 3707 17436
rect 3707 17380 3711 17436
rect 3647 17376 3711 17380
rect 3727 17436 3791 17440
rect 3727 17380 3731 17436
rect 3731 17380 3787 17436
rect 3787 17380 3791 17436
rect 3727 17376 3791 17380
rect 3807 17436 3871 17440
rect 3807 17380 3811 17436
rect 3811 17380 3867 17436
rect 3867 17380 3871 17436
rect 3807 17376 3871 17380
rect 3887 17436 3951 17440
rect 3887 17380 3891 17436
rect 3891 17380 3947 17436
rect 3947 17380 3951 17436
rect 3887 17376 3951 17380
rect 7718 17436 7782 17440
rect 7718 17380 7722 17436
rect 7722 17380 7778 17436
rect 7778 17380 7782 17436
rect 7718 17376 7782 17380
rect 7798 17436 7862 17440
rect 7798 17380 7802 17436
rect 7802 17380 7858 17436
rect 7858 17380 7862 17436
rect 7798 17376 7862 17380
rect 7878 17436 7942 17440
rect 7878 17380 7882 17436
rect 7882 17380 7938 17436
rect 7938 17380 7942 17436
rect 7878 17376 7942 17380
rect 7958 17436 8022 17440
rect 7958 17380 7962 17436
rect 7962 17380 8018 17436
rect 8018 17380 8022 17436
rect 7958 17376 8022 17380
rect 11789 17436 11853 17440
rect 11789 17380 11793 17436
rect 11793 17380 11849 17436
rect 11849 17380 11853 17436
rect 11789 17376 11853 17380
rect 11869 17436 11933 17440
rect 11869 17380 11873 17436
rect 11873 17380 11929 17436
rect 11929 17380 11933 17436
rect 11869 17376 11933 17380
rect 11949 17436 12013 17440
rect 11949 17380 11953 17436
rect 11953 17380 12009 17436
rect 12009 17380 12013 17436
rect 11949 17376 12013 17380
rect 12029 17436 12093 17440
rect 12029 17380 12033 17436
rect 12033 17380 12089 17436
rect 12089 17380 12093 17436
rect 12029 17376 12093 17380
rect 15860 17436 15924 17440
rect 15860 17380 15864 17436
rect 15864 17380 15920 17436
rect 15920 17380 15924 17436
rect 15860 17376 15924 17380
rect 15940 17436 16004 17440
rect 15940 17380 15944 17436
rect 15944 17380 16000 17436
rect 16000 17380 16004 17436
rect 15940 17376 16004 17380
rect 16020 17436 16084 17440
rect 16020 17380 16024 17436
rect 16024 17380 16080 17436
rect 16080 17380 16084 17436
rect 16020 17376 16084 17380
rect 16100 17436 16164 17440
rect 16100 17380 16104 17436
rect 16104 17380 16160 17436
rect 16160 17380 16164 17436
rect 16100 17376 16164 17380
rect 2987 16892 3051 16896
rect 2987 16836 2991 16892
rect 2991 16836 3047 16892
rect 3047 16836 3051 16892
rect 2987 16832 3051 16836
rect 3067 16892 3131 16896
rect 3067 16836 3071 16892
rect 3071 16836 3127 16892
rect 3127 16836 3131 16892
rect 3067 16832 3131 16836
rect 3147 16892 3211 16896
rect 3147 16836 3151 16892
rect 3151 16836 3207 16892
rect 3207 16836 3211 16892
rect 3147 16832 3211 16836
rect 3227 16892 3291 16896
rect 3227 16836 3231 16892
rect 3231 16836 3287 16892
rect 3287 16836 3291 16892
rect 3227 16832 3291 16836
rect 7058 16892 7122 16896
rect 7058 16836 7062 16892
rect 7062 16836 7118 16892
rect 7118 16836 7122 16892
rect 7058 16832 7122 16836
rect 7138 16892 7202 16896
rect 7138 16836 7142 16892
rect 7142 16836 7198 16892
rect 7198 16836 7202 16892
rect 7138 16832 7202 16836
rect 7218 16892 7282 16896
rect 7218 16836 7222 16892
rect 7222 16836 7278 16892
rect 7278 16836 7282 16892
rect 7218 16832 7282 16836
rect 7298 16892 7362 16896
rect 7298 16836 7302 16892
rect 7302 16836 7358 16892
rect 7358 16836 7362 16892
rect 7298 16832 7362 16836
rect 11129 16892 11193 16896
rect 11129 16836 11133 16892
rect 11133 16836 11189 16892
rect 11189 16836 11193 16892
rect 11129 16832 11193 16836
rect 11209 16892 11273 16896
rect 11209 16836 11213 16892
rect 11213 16836 11269 16892
rect 11269 16836 11273 16892
rect 11209 16832 11273 16836
rect 11289 16892 11353 16896
rect 11289 16836 11293 16892
rect 11293 16836 11349 16892
rect 11349 16836 11353 16892
rect 11289 16832 11353 16836
rect 11369 16892 11433 16896
rect 11369 16836 11373 16892
rect 11373 16836 11429 16892
rect 11429 16836 11433 16892
rect 11369 16832 11433 16836
rect 15200 16892 15264 16896
rect 15200 16836 15204 16892
rect 15204 16836 15260 16892
rect 15260 16836 15264 16892
rect 15200 16832 15264 16836
rect 15280 16892 15344 16896
rect 15280 16836 15284 16892
rect 15284 16836 15340 16892
rect 15340 16836 15344 16892
rect 15280 16832 15344 16836
rect 15360 16892 15424 16896
rect 15360 16836 15364 16892
rect 15364 16836 15420 16892
rect 15420 16836 15424 16892
rect 15360 16832 15424 16836
rect 15440 16892 15504 16896
rect 15440 16836 15444 16892
rect 15444 16836 15500 16892
rect 15500 16836 15504 16892
rect 15440 16832 15504 16836
rect 3647 16348 3711 16352
rect 3647 16292 3651 16348
rect 3651 16292 3707 16348
rect 3707 16292 3711 16348
rect 3647 16288 3711 16292
rect 3727 16348 3791 16352
rect 3727 16292 3731 16348
rect 3731 16292 3787 16348
rect 3787 16292 3791 16348
rect 3727 16288 3791 16292
rect 3807 16348 3871 16352
rect 3807 16292 3811 16348
rect 3811 16292 3867 16348
rect 3867 16292 3871 16348
rect 3807 16288 3871 16292
rect 3887 16348 3951 16352
rect 3887 16292 3891 16348
rect 3891 16292 3947 16348
rect 3947 16292 3951 16348
rect 3887 16288 3951 16292
rect 7718 16348 7782 16352
rect 7718 16292 7722 16348
rect 7722 16292 7778 16348
rect 7778 16292 7782 16348
rect 7718 16288 7782 16292
rect 7798 16348 7862 16352
rect 7798 16292 7802 16348
rect 7802 16292 7858 16348
rect 7858 16292 7862 16348
rect 7798 16288 7862 16292
rect 7878 16348 7942 16352
rect 7878 16292 7882 16348
rect 7882 16292 7938 16348
rect 7938 16292 7942 16348
rect 7878 16288 7942 16292
rect 7958 16348 8022 16352
rect 7958 16292 7962 16348
rect 7962 16292 8018 16348
rect 8018 16292 8022 16348
rect 7958 16288 8022 16292
rect 11789 16348 11853 16352
rect 11789 16292 11793 16348
rect 11793 16292 11849 16348
rect 11849 16292 11853 16348
rect 11789 16288 11853 16292
rect 11869 16348 11933 16352
rect 11869 16292 11873 16348
rect 11873 16292 11929 16348
rect 11929 16292 11933 16348
rect 11869 16288 11933 16292
rect 11949 16348 12013 16352
rect 11949 16292 11953 16348
rect 11953 16292 12009 16348
rect 12009 16292 12013 16348
rect 11949 16288 12013 16292
rect 12029 16348 12093 16352
rect 12029 16292 12033 16348
rect 12033 16292 12089 16348
rect 12089 16292 12093 16348
rect 12029 16288 12093 16292
rect 15860 16348 15924 16352
rect 15860 16292 15864 16348
rect 15864 16292 15920 16348
rect 15920 16292 15924 16348
rect 15860 16288 15924 16292
rect 15940 16348 16004 16352
rect 15940 16292 15944 16348
rect 15944 16292 16000 16348
rect 16000 16292 16004 16348
rect 15940 16288 16004 16292
rect 16020 16348 16084 16352
rect 16020 16292 16024 16348
rect 16024 16292 16080 16348
rect 16080 16292 16084 16348
rect 16020 16288 16084 16292
rect 16100 16348 16164 16352
rect 16100 16292 16104 16348
rect 16104 16292 16160 16348
rect 16160 16292 16164 16348
rect 16100 16288 16164 16292
rect 2987 15804 3051 15808
rect 2987 15748 2991 15804
rect 2991 15748 3047 15804
rect 3047 15748 3051 15804
rect 2987 15744 3051 15748
rect 3067 15804 3131 15808
rect 3067 15748 3071 15804
rect 3071 15748 3127 15804
rect 3127 15748 3131 15804
rect 3067 15744 3131 15748
rect 3147 15804 3211 15808
rect 3147 15748 3151 15804
rect 3151 15748 3207 15804
rect 3207 15748 3211 15804
rect 3147 15744 3211 15748
rect 3227 15804 3291 15808
rect 3227 15748 3231 15804
rect 3231 15748 3287 15804
rect 3287 15748 3291 15804
rect 3227 15744 3291 15748
rect 7058 15804 7122 15808
rect 7058 15748 7062 15804
rect 7062 15748 7118 15804
rect 7118 15748 7122 15804
rect 7058 15744 7122 15748
rect 7138 15804 7202 15808
rect 7138 15748 7142 15804
rect 7142 15748 7198 15804
rect 7198 15748 7202 15804
rect 7138 15744 7202 15748
rect 7218 15804 7282 15808
rect 7218 15748 7222 15804
rect 7222 15748 7278 15804
rect 7278 15748 7282 15804
rect 7218 15744 7282 15748
rect 7298 15804 7362 15808
rect 7298 15748 7302 15804
rect 7302 15748 7358 15804
rect 7358 15748 7362 15804
rect 7298 15744 7362 15748
rect 11129 15804 11193 15808
rect 11129 15748 11133 15804
rect 11133 15748 11189 15804
rect 11189 15748 11193 15804
rect 11129 15744 11193 15748
rect 11209 15804 11273 15808
rect 11209 15748 11213 15804
rect 11213 15748 11269 15804
rect 11269 15748 11273 15804
rect 11209 15744 11273 15748
rect 11289 15804 11353 15808
rect 11289 15748 11293 15804
rect 11293 15748 11349 15804
rect 11349 15748 11353 15804
rect 11289 15744 11353 15748
rect 11369 15804 11433 15808
rect 11369 15748 11373 15804
rect 11373 15748 11429 15804
rect 11429 15748 11433 15804
rect 11369 15744 11433 15748
rect 15200 15804 15264 15808
rect 15200 15748 15204 15804
rect 15204 15748 15260 15804
rect 15260 15748 15264 15804
rect 15200 15744 15264 15748
rect 15280 15804 15344 15808
rect 15280 15748 15284 15804
rect 15284 15748 15340 15804
rect 15340 15748 15344 15804
rect 15280 15744 15344 15748
rect 15360 15804 15424 15808
rect 15360 15748 15364 15804
rect 15364 15748 15420 15804
rect 15420 15748 15424 15804
rect 15360 15744 15424 15748
rect 15440 15804 15504 15808
rect 15440 15748 15444 15804
rect 15444 15748 15500 15804
rect 15500 15748 15504 15804
rect 15440 15744 15504 15748
rect 3647 15260 3711 15264
rect 3647 15204 3651 15260
rect 3651 15204 3707 15260
rect 3707 15204 3711 15260
rect 3647 15200 3711 15204
rect 3727 15260 3791 15264
rect 3727 15204 3731 15260
rect 3731 15204 3787 15260
rect 3787 15204 3791 15260
rect 3727 15200 3791 15204
rect 3807 15260 3871 15264
rect 3807 15204 3811 15260
rect 3811 15204 3867 15260
rect 3867 15204 3871 15260
rect 3807 15200 3871 15204
rect 3887 15260 3951 15264
rect 3887 15204 3891 15260
rect 3891 15204 3947 15260
rect 3947 15204 3951 15260
rect 3887 15200 3951 15204
rect 7718 15260 7782 15264
rect 7718 15204 7722 15260
rect 7722 15204 7778 15260
rect 7778 15204 7782 15260
rect 7718 15200 7782 15204
rect 7798 15260 7862 15264
rect 7798 15204 7802 15260
rect 7802 15204 7858 15260
rect 7858 15204 7862 15260
rect 7798 15200 7862 15204
rect 7878 15260 7942 15264
rect 7878 15204 7882 15260
rect 7882 15204 7938 15260
rect 7938 15204 7942 15260
rect 7878 15200 7942 15204
rect 7958 15260 8022 15264
rect 7958 15204 7962 15260
rect 7962 15204 8018 15260
rect 8018 15204 8022 15260
rect 7958 15200 8022 15204
rect 11789 15260 11853 15264
rect 11789 15204 11793 15260
rect 11793 15204 11849 15260
rect 11849 15204 11853 15260
rect 11789 15200 11853 15204
rect 11869 15260 11933 15264
rect 11869 15204 11873 15260
rect 11873 15204 11929 15260
rect 11929 15204 11933 15260
rect 11869 15200 11933 15204
rect 11949 15260 12013 15264
rect 11949 15204 11953 15260
rect 11953 15204 12009 15260
rect 12009 15204 12013 15260
rect 11949 15200 12013 15204
rect 12029 15260 12093 15264
rect 12029 15204 12033 15260
rect 12033 15204 12089 15260
rect 12089 15204 12093 15260
rect 12029 15200 12093 15204
rect 15860 15260 15924 15264
rect 15860 15204 15864 15260
rect 15864 15204 15920 15260
rect 15920 15204 15924 15260
rect 15860 15200 15924 15204
rect 15940 15260 16004 15264
rect 15940 15204 15944 15260
rect 15944 15204 16000 15260
rect 16000 15204 16004 15260
rect 15940 15200 16004 15204
rect 16020 15260 16084 15264
rect 16020 15204 16024 15260
rect 16024 15204 16080 15260
rect 16080 15204 16084 15260
rect 16020 15200 16084 15204
rect 16100 15260 16164 15264
rect 16100 15204 16104 15260
rect 16104 15204 16160 15260
rect 16160 15204 16164 15260
rect 16100 15200 16164 15204
rect 2987 14716 3051 14720
rect 2987 14660 2991 14716
rect 2991 14660 3047 14716
rect 3047 14660 3051 14716
rect 2987 14656 3051 14660
rect 3067 14716 3131 14720
rect 3067 14660 3071 14716
rect 3071 14660 3127 14716
rect 3127 14660 3131 14716
rect 3067 14656 3131 14660
rect 3147 14716 3211 14720
rect 3147 14660 3151 14716
rect 3151 14660 3207 14716
rect 3207 14660 3211 14716
rect 3147 14656 3211 14660
rect 3227 14716 3291 14720
rect 3227 14660 3231 14716
rect 3231 14660 3287 14716
rect 3287 14660 3291 14716
rect 3227 14656 3291 14660
rect 7058 14716 7122 14720
rect 7058 14660 7062 14716
rect 7062 14660 7118 14716
rect 7118 14660 7122 14716
rect 7058 14656 7122 14660
rect 7138 14716 7202 14720
rect 7138 14660 7142 14716
rect 7142 14660 7198 14716
rect 7198 14660 7202 14716
rect 7138 14656 7202 14660
rect 7218 14716 7282 14720
rect 7218 14660 7222 14716
rect 7222 14660 7278 14716
rect 7278 14660 7282 14716
rect 7218 14656 7282 14660
rect 7298 14716 7362 14720
rect 7298 14660 7302 14716
rect 7302 14660 7358 14716
rect 7358 14660 7362 14716
rect 7298 14656 7362 14660
rect 11129 14716 11193 14720
rect 11129 14660 11133 14716
rect 11133 14660 11189 14716
rect 11189 14660 11193 14716
rect 11129 14656 11193 14660
rect 11209 14716 11273 14720
rect 11209 14660 11213 14716
rect 11213 14660 11269 14716
rect 11269 14660 11273 14716
rect 11209 14656 11273 14660
rect 11289 14716 11353 14720
rect 11289 14660 11293 14716
rect 11293 14660 11349 14716
rect 11349 14660 11353 14716
rect 11289 14656 11353 14660
rect 11369 14716 11433 14720
rect 11369 14660 11373 14716
rect 11373 14660 11429 14716
rect 11429 14660 11433 14716
rect 11369 14656 11433 14660
rect 15200 14716 15264 14720
rect 15200 14660 15204 14716
rect 15204 14660 15260 14716
rect 15260 14660 15264 14716
rect 15200 14656 15264 14660
rect 15280 14716 15344 14720
rect 15280 14660 15284 14716
rect 15284 14660 15340 14716
rect 15340 14660 15344 14716
rect 15280 14656 15344 14660
rect 15360 14716 15424 14720
rect 15360 14660 15364 14716
rect 15364 14660 15420 14716
rect 15420 14660 15424 14716
rect 15360 14656 15424 14660
rect 15440 14716 15504 14720
rect 15440 14660 15444 14716
rect 15444 14660 15500 14716
rect 15500 14660 15504 14716
rect 15440 14656 15504 14660
rect 3647 14172 3711 14176
rect 3647 14116 3651 14172
rect 3651 14116 3707 14172
rect 3707 14116 3711 14172
rect 3647 14112 3711 14116
rect 3727 14172 3791 14176
rect 3727 14116 3731 14172
rect 3731 14116 3787 14172
rect 3787 14116 3791 14172
rect 3727 14112 3791 14116
rect 3807 14172 3871 14176
rect 3807 14116 3811 14172
rect 3811 14116 3867 14172
rect 3867 14116 3871 14172
rect 3807 14112 3871 14116
rect 3887 14172 3951 14176
rect 3887 14116 3891 14172
rect 3891 14116 3947 14172
rect 3947 14116 3951 14172
rect 3887 14112 3951 14116
rect 7718 14172 7782 14176
rect 7718 14116 7722 14172
rect 7722 14116 7778 14172
rect 7778 14116 7782 14172
rect 7718 14112 7782 14116
rect 7798 14172 7862 14176
rect 7798 14116 7802 14172
rect 7802 14116 7858 14172
rect 7858 14116 7862 14172
rect 7798 14112 7862 14116
rect 7878 14172 7942 14176
rect 7878 14116 7882 14172
rect 7882 14116 7938 14172
rect 7938 14116 7942 14172
rect 7878 14112 7942 14116
rect 7958 14172 8022 14176
rect 7958 14116 7962 14172
rect 7962 14116 8018 14172
rect 8018 14116 8022 14172
rect 7958 14112 8022 14116
rect 11789 14172 11853 14176
rect 11789 14116 11793 14172
rect 11793 14116 11849 14172
rect 11849 14116 11853 14172
rect 11789 14112 11853 14116
rect 11869 14172 11933 14176
rect 11869 14116 11873 14172
rect 11873 14116 11929 14172
rect 11929 14116 11933 14172
rect 11869 14112 11933 14116
rect 11949 14172 12013 14176
rect 11949 14116 11953 14172
rect 11953 14116 12009 14172
rect 12009 14116 12013 14172
rect 11949 14112 12013 14116
rect 12029 14172 12093 14176
rect 12029 14116 12033 14172
rect 12033 14116 12089 14172
rect 12089 14116 12093 14172
rect 12029 14112 12093 14116
rect 15860 14172 15924 14176
rect 15860 14116 15864 14172
rect 15864 14116 15920 14172
rect 15920 14116 15924 14172
rect 15860 14112 15924 14116
rect 15940 14172 16004 14176
rect 15940 14116 15944 14172
rect 15944 14116 16000 14172
rect 16000 14116 16004 14172
rect 15940 14112 16004 14116
rect 16020 14172 16084 14176
rect 16020 14116 16024 14172
rect 16024 14116 16080 14172
rect 16080 14116 16084 14172
rect 16020 14112 16084 14116
rect 16100 14172 16164 14176
rect 16100 14116 16104 14172
rect 16104 14116 16160 14172
rect 16160 14116 16164 14172
rect 16100 14112 16164 14116
rect 2987 13628 3051 13632
rect 2987 13572 2991 13628
rect 2991 13572 3047 13628
rect 3047 13572 3051 13628
rect 2987 13568 3051 13572
rect 3067 13628 3131 13632
rect 3067 13572 3071 13628
rect 3071 13572 3127 13628
rect 3127 13572 3131 13628
rect 3067 13568 3131 13572
rect 3147 13628 3211 13632
rect 3147 13572 3151 13628
rect 3151 13572 3207 13628
rect 3207 13572 3211 13628
rect 3147 13568 3211 13572
rect 3227 13628 3291 13632
rect 3227 13572 3231 13628
rect 3231 13572 3287 13628
rect 3287 13572 3291 13628
rect 3227 13568 3291 13572
rect 7058 13628 7122 13632
rect 7058 13572 7062 13628
rect 7062 13572 7118 13628
rect 7118 13572 7122 13628
rect 7058 13568 7122 13572
rect 7138 13628 7202 13632
rect 7138 13572 7142 13628
rect 7142 13572 7198 13628
rect 7198 13572 7202 13628
rect 7138 13568 7202 13572
rect 7218 13628 7282 13632
rect 7218 13572 7222 13628
rect 7222 13572 7278 13628
rect 7278 13572 7282 13628
rect 7218 13568 7282 13572
rect 7298 13628 7362 13632
rect 7298 13572 7302 13628
rect 7302 13572 7358 13628
rect 7358 13572 7362 13628
rect 7298 13568 7362 13572
rect 11129 13628 11193 13632
rect 11129 13572 11133 13628
rect 11133 13572 11189 13628
rect 11189 13572 11193 13628
rect 11129 13568 11193 13572
rect 11209 13628 11273 13632
rect 11209 13572 11213 13628
rect 11213 13572 11269 13628
rect 11269 13572 11273 13628
rect 11209 13568 11273 13572
rect 11289 13628 11353 13632
rect 11289 13572 11293 13628
rect 11293 13572 11349 13628
rect 11349 13572 11353 13628
rect 11289 13568 11353 13572
rect 11369 13628 11433 13632
rect 11369 13572 11373 13628
rect 11373 13572 11429 13628
rect 11429 13572 11433 13628
rect 11369 13568 11433 13572
rect 15200 13628 15264 13632
rect 15200 13572 15204 13628
rect 15204 13572 15260 13628
rect 15260 13572 15264 13628
rect 15200 13568 15264 13572
rect 15280 13628 15344 13632
rect 15280 13572 15284 13628
rect 15284 13572 15340 13628
rect 15340 13572 15344 13628
rect 15280 13568 15344 13572
rect 15360 13628 15424 13632
rect 15360 13572 15364 13628
rect 15364 13572 15420 13628
rect 15420 13572 15424 13628
rect 15360 13568 15424 13572
rect 15440 13628 15504 13632
rect 15440 13572 15444 13628
rect 15444 13572 15500 13628
rect 15500 13572 15504 13628
rect 15440 13568 15504 13572
rect 3647 13084 3711 13088
rect 3647 13028 3651 13084
rect 3651 13028 3707 13084
rect 3707 13028 3711 13084
rect 3647 13024 3711 13028
rect 3727 13084 3791 13088
rect 3727 13028 3731 13084
rect 3731 13028 3787 13084
rect 3787 13028 3791 13084
rect 3727 13024 3791 13028
rect 3807 13084 3871 13088
rect 3807 13028 3811 13084
rect 3811 13028 3867 13084
rect 3867 13028 3871 13084
rect 3807 13024 3871 13028
rect 3887 13084 3951 13088
rect 3887 13028 3891 13084
rect 3891 13028 3947 13084
rect 3947 13028 3951 13084
rect 3887 13024 3951 13028
rect 7718 13084 7782 13088
rect 7718 13028 7722 13084
rect 7722 13028 7778 13084
rect 7778 13028 7782 13084
rect 7718 13024 7782 13028
rect 7798 13084 7862 13088
rect 7798 13028 7802 13084
rect 7802 13028 7858 13084
rect 7858 13028 7862 13084
rect 7798 13024 7862 13028
rect 7878 13084 7942 13088
rect 7878 13028 7882 13084
rect 7882 13028 7938 13084
rect 7938 13028 7942 13084
rect 7878 13024 7942 13028
rect 7958 13084 8022 13088
rect 7958 13028 7962 13084
rect 7962 13028 8018 13084
rect 8018 13028 8022 13084
rect 7958 13024 8022 13028
rect 11789 13084 11853 13088
rect 11789 13028 11793 13084
rect 11793 13028 11849 13084
rect 11849 13028 11853 13084
rect 11789 13024 11853 13028
rect 11869 13084 11933 13088
rect 11869 13028 11873 13084
rect 11873 13028 11929 13084
rect 11929 13028 11933 13084
rect 11869 13024 11933 13028
rect 11949 13084 12013 13088
rect 11949 13028 11953 13084
rect 11953 13028 12009 13084
rect 12009 13028 12013 13084
rect 11949 13024 12013 13028
rect 12029 13084 12093 13088
rect 12029 13028 12033 13084
rect 12033 13028 12089 13084
rect 12089 13028 12093 13084
rect 12029 13024 12093 13028
rect 15860 13084 15924 13088
rect 15860 13028 15864 13084
rect 15864 13028 15920 13084
rect 15920 13028 15924 13084
rect 15860 13024 15924 13028
rect 15940 13084 16004 13088
rect 15940 13028 15944 13084
rect 15944 13028 16000 13084
rect 16000 13028 16004 13084
rect 15940 13024 16004 13028
rect 16020 13084 16084 13088
rect 16020 13028 16024 13084
rect 16024 13028 16080 13084
rect 16080 13028 16084 13084
rect 16020 13024 16084 13028
rect 16100 13084 16164 13088
rect 16100 13028 16104 13084
rect 16104 13028 16160 13084
rect 16160 13028 16164 13084
rect 16100 13024 16164 13028
rect 2987 12540 3051 12544
rect 2987 12484 2991 12540
rect 2991 12484 3047 12540
rect 3047 12484 3051 12540
rect 2987 12480 3051 12484
rect 3067 12540 3131 12544
rect 3067 12484 3071 12540
rect 3071 12484 3127 12540
rect 3127 12484 3131 12540
rect 3067 12480 3131 12484
rect 3147 12540 3211 12544
rect 3147 12484 3151 12540
rect 3151 12484 3207 12540
rect 3207 12484 3211 12540
rect 3147 12480 3211 12484
rect 3227 12540 3291 12544
rect 3227 12484 3231 12540
rect 3231 12484 3287 12540
rect 3287 12484 3291 12540
rect 3227 12480 3291 12484
rect 7058 12540 7122 12544
rect 7058 12484 7062 12540
rect 7062 12484 7118 12540
rect 7118 12484 7122 12540
rect 7058 12480 7122 12484
rect 7138 12540 7202 12544
rect 7138 12484 7142 12540
rect 7142 12484 7198 12540
rect 7198 12484 7202 12540
rect 7138 12480 7202 12484
rect 7218 12540 7282 12544
rect 7218 12484 7222 12540
rect 7222 12484 7278 12540
rect 7278 12484 7282 12540
rect 7218 12480 7282 12484
rect 7298 12540 7362 12544
rect 7298 12484 7302 12540
rect 7302 12484 7358 12540
rect 7358 12484 7362 12540
rect 7298 12480 7362 12484
rect 11129 12540 11193 12544
rect 11129 12484 11133 12540
rect 11133 12484 11189 12540
rect 11189 12484 11193 12540
rect 11129 12480 11193 12484
rect 11209 12540 11273 12544
rect 11209 12484 11213 12540
rect 11213 12484 11269 12540
rect 11269 12484 11273 12540
rect 11209 12480 11273 12484
rect 11289 12540 11353 12544
rect 11289 12484 11293 12540
rect 11293 12484 11349 12540
rect 11349 12484 11353 12540
rect 11289 12480 11353 12484
rect 11369 12540 11433 12544
rect 11369 12484 11373 12540
rect 11373 12484 11429 12540
rect 11429 12484 11433 12540
rect 11369 12480 11433 12484
rect 15200 12540 15264 12544
rect 15200 12484 15204 12540
rect 15204 12484 15260 12540
rect 15260 12484 15264 12540
rect 15200 12480 15264 12484
rect 15280 12540 15344 12544
rect 15280 12484 15284 12540
rect 15284 12484 15340 12540
rect 15340 12484 15344 12540
rect 15280 12480 15344 12484
rect 15360 12540 15424 12544
rect 15360 12484 15364 12540
rect 15364 12484 15420 12540
rect 15420 12484 15424 12540
rect 15360 12480 15424 12484
rect 15440 12540 15504 12544
rect 15440 12484 15444 12540
rect 15444 12484 15500 12540
rect 15500 12484 15504 12540
rect 15440 12480 15504 12484
rect 3647 11996 3711 12000
rect 3647 11940 3651 11996
rect 3651 11940 3707 11996
rect 3707 11940 3711 11996
rect 3647 11936 3711 11940
rect 3727 11996 3791 12000
rect 3727 11940 3731 11996
rect 3731 11940 3787 11996
rect 3787 11940 3791 11996
rect 3727 11936 3791 11940
rect 3807 11996 3871 12000
rect 3807 11940 3811 11996
rect 3811 11940 3867 11996
rect 3867 11940 3871 11996
rect 3807 11936 3871 11940
rect 3887 11996 3951 12000
rect 3887 11940 3891 11996
rect 3891 11940 3947 11996
rect 3947 11940 3951 11996
rect 3887 11936 3951 11940
rect 7718 11996 7782 12000
rect 7718 11940 7722 11996
rect 7722 11940 7778 11996
rect 7778 11940 7782 11996
rect 7718 11936 7782 11940
rect 7798 11996 7862 12000
rect 7798 11940 7802 11996
rect 7802 11940 7858 11996
rect 7858 11940 7862 11996
rect 7798 11936 7862 11940
rect 7878 11996 7942 12000
rect 7878 11940 7882 11996
rect 7882 11940 7938 11996
rect 7938 11940 7942 11996
rect 7878 11936 7942 11940
rect 7958 11996 8022 12000
rect 7958 11940 7962 11996
rect 7962 11940 8018 11996
rect 8018 11940 8022 11996
rect 7958 11936 8022 11940
rect 11789 11996 11853 12000
rect 11789 11940 11793 11996
rect 11793 11940 11849 11996
rect 11849 11940 11853 11996
rect 11789 11936 11853 11940
rect 11869 11996 11933 12000
rect 11869 11940 11873 11996
rect 11873 11940 11929 11996
rect 11929 11940 11933 11996
rect 11869 11936 11933 11940
rect 11949 11996 12013 12000
rect 11949 11940 11953 11996
rect 11953 11940 12009 11996
rect 12009 11940 12013 11996
rect 11949 11936 12013 11940
rect 12029 11996 12093 12000
rect 12029 11940 12033 11996
rect 12033 11940 12089 11996
rect 12089 11940 12093 11996
rect 12029 11936 12093 11940
rect 15860 11996 15924 12000
rect 15860 11940 15864 11996
rect 15864 11940 15920 11996
rect 15920 11940 15924 11996
rect 15860 11936 15924 11940
rect 15940 11996 16004 12000
rect 15940 11940 15944 11996
rect 15944 11940 16000 11996
rect 16000 11940 16004 11996
rect 15940 11936 16004 11940
rect 16020 11996 16084 12000
rect 16020 11940 16024 11996
rect 16024 11940 16080 11996
rect 16080 11940 16084 11996
rect 16020 11936 16084 11940
rect 16100 11996 16164 12000
rect 16100 11940 16104 11996
rect 16104 11940 16160 11996
rect 16160 11940 16164 11996
rect 16100 11936 16164 11940
rect 2987 11452 3051 11456
rect 2987 11396 2991 11452
rect 2991 11396 3047 11452
rect 3047 11396 3051 11452
rect 2987 11392 3051 11396
rect 3067 11452 3131 11456
rect 3067 11396 3071 11452
rect 3071 11396 3127 11452
rect 3127 11396 3131 11452
rect 3067 11392 3131 11396
rect 3147 11452 3211 11456
rect 3147 11396 3151 11452
rect 3151 11396 3207 11452
rect 3207 11396 3211 11452
rect 3147 11392 3211 11396
rect 3227 11452 3291 11456
rect 3227 11396 3231 11452
rect 3231 11396 3287 11452
rect 3287 11396 3291 11452
rect 3227 11392 3291 11396
rect 7058 11452 7122 11456
rect 7058 11396 7062 11452
rect 7062 11396 7118 11452
rect 7118 11396 7122 11452
rect 7058 11392 7122 11396
rect 7138 11452 7202 11456
rect 7138 11396 7142 11452
rect 7142 11396 7198 11452
rect 7198 11396 7202 11452
rect 7138 11392 7202 11396
rect 7218 11452 7282 11456
rect 7218 11396 7222 11452
rect 7222 11396 7278 11452
rect 7278 11396 7282 11452
rect 7218 11392 7282 11396
rect 7298 11452 7362 11456
rect 7298 11396 7302 11452
rect 7302 11396 7358 11452
rect 7358 11396 7362 11452
rect 7298 11392 7362 11396
rect 11129 11452 11193 11456
rect 11129 11396 11133 11452
rect 11133 11396 11189 11452
rect 11189 11396 11193 11452
rect 11129 11392 11193 11396
rect 11209 11452 11273 11456
rect 11209 11396 11213 11452
rect 11213 11396 11269 11452
rect 11269 11396 11273 11452
rect 11209 11392 11273 11396
rect 11289 11452 11353 11456
rect 11289 11396 11293 11452
rect 11293 11396 11349 11452
rect 11349 11396 11353 11452
rect 11289 11392 11353 11396
rect 11369 11452 11433 11456
rect 11369 11396 11373 11452
rect 11373 11396 11429 11452
rect 11429 11396 11433 11452
rect 11369 11392 11433 11396
rect 15200 11452 15264 11456
rect 15200 11396 15204 11452
rect 15204 11396 15260 11452
rect 15260 11396 15264 11452
rect 15200 11392 15264 11396
rect 15280 11452 15344 11456
rect 15280 11396 15284 11452
rect 15284 11396 15340 11452
rect 15340 11396 15344 11452
rect 15280 11392 15344 11396
rect 15360 11452 15424 11456
rect 15360 11396 15364 11452
rect 15364 11396 15420 11452
rect 15420 11396 15424 11452
rect 15360 11392 15424 11396
rect 15440 11452 15504 11456
rect 15440 11396 15444 11452
rect 15444 11396 15500 11452
rect 15500 11396 15504 11452
rect 15440 11392 15504 11396
rect 3647 10908 3711 10912
rect 3647 10852 3651 10908
rect 3651 10852 3707 10908
rect 3707 10852 3711 10908
rect 3647 10848 3711 10852
rect 3727 10908 3791 10912
rect 3727 10852 3731 10908
rect 3731 10852 3787 10908
rect 3787 10852 3791 10908
rect 3727 10848 3791 10852
rect 3807 10908 3871 10912
rect 3807 10852 3811 10908
rect 3811 10852 3867 10908
rect 3867 10852 3871 10908
rect 3807 10848 3871 10852
rect 3887 10908 3951 10912
rect 3887 10852 3891 10908
rect 3891 10852 3947 10908
rect 3947 10852 3951 10908
rect 3887 10848 3951 10852
rect 7718 10908 7782 10912
rect 7718 10852 7722 10908
rect 7722 10852 7778 10908
rect 7778 10852 7782 10908
rect 7718 10848 7782 10852
rect 7798 10908 7862 10912
rect 7798 10852 7802 10908
rect 7802 10852 7858 10908
rect 7858 10852 7862 10908
rect 7798 10848 7862 10852
rect 7878 10908 7942 10912
rect 7878 10852 7882 10908
rect 7882 10852 7938 10908
rect 7938 10852 7942 10908
rect 7878 10848 7942 10852
rect 7958 10908 8022 10912
rect 7958 10852 7962 10908
rect 7962 10852 8018 10908
rect 8018 10852 8022 10908
rect 7958 10848 8022 10852
rect 11789 10908 11853 10912
rect 11789 10852 11793 10908
rect 11793 10852 11849 10908
rect 11849 10852 11853 10908
rect 11789 10848 11853 10852
rect 11869 10908 11933 10912
rect 11869 10852 11873 10908
rect 11873 10852 11929 10908
rect 11929 10852 11933 10908
rect 11869 10848 11933 10852
rect 11949 10908 12013 10912
rect 11949 10852 11953 10908
rect 11953 10852 12009 10908
rect 12009 10852 12013 10908
rect 11949 10848 12013 10852
rect 12029 10908 12093 10912
rect 12029 10852 12033 10908
rect 12033 10852 12089 10908
rect 12089 10852 12093 10908
rect 12029 10848 12093 10852
rect 15860 10908 15924 10912
rect 15860 10852 15864 10908
rect 15864 10852 15920 10908
rect 15920 10852 15924 10908
rect 15860 10848 15924 10852
rect 15940 10908 16004 10912
rect 15940 10852 15944 10908
rect 15944 10852 16000 10908
rect 16000 10852 16004 10908
rect 15940 10848 16004 10852
rect 16020 10908 16084 10912
rect 16020 10852 16024 10908
rect 16024 10852 16080 10908
rect 16080 10852 16084 10908
rect 16020 10848 16084 10852
rect 16100 10908 16164 10912
rect 16100 10852 16104 10908
rect 16104 10852 16160 10908
rect 16160 10852 16164 10908
rect 16100 10848 16164 10852
rect 2987 10364 3051 10368
rect 2987 10308 2991 10364
rect 2991 10308 3047 10364
rect 3047 10308 3051 10364
rect 2987 10304 3051 10308
rect 3067 10364 3131 10368
rect 3067 10308 3071 10364
rect 3071 10308 3127 10364
rect 3127 10308 3131 10364
rect 3067 10304 3131 10308
rect 3147 10364 3211 10368
rect 3147 10308 3151 10364
rect 3151 10308 3207 10364
rect 3207 10308 3211 10364
rect 3147 10304 3211 10308
rect 3227 10364 3291 10368
rect 3227 10308 3231 10364
rect 3231 10308 3287 10364
rect 3287 10308 3291 10364
rect 3227 10304 3291 10308
rect 7058 10364 7122 10368
rect 7058 10308 7062 10364
rect 7062 10308 7118 10364
rect 7118 10308 7122 10364
rect 7058 10304 7122 10308
rect 7138 10364 7202 10368
rect 7138 10308 7142 10364
rect 7142 10308 7198 10364
rect 7198 10308 7202 10364
rect 7138 10304 7202 10308
rect 7218 10364 7282 10368
rect 7218 10308 7222 10364
rect 7222 10308 7278 10364
rect 7278 10308 7282 10364
rect 7218 10304 7282 10308
rect 7298 10364 7362 10368
rect 7298 10308 7302 10364
rect 7302 10308 7358 10364
rect 7358 10308 7362 10364
rect 7298 10304 7362 10308
rect 11129 10364 11193 10368
rect 11129 10308 11133 10364
rect 11133 10308 11189 10364
rect 11189 10308 11193 10364
rect 11129 10304 11193 10308
rect 11209 10364 11273 10368
rect 11209 10308 11213 10364
rect 11213 10308 11269 10364
rect 11269 10308 11273 10364
rect 11209 10304 11273 10308
rect 11289 10364 11353 10368
rect 11289 10308 11293 10364
rect 11293 10308 11349 10364
rect 11349 10308 11353 10364
rect 11289 10304 11353 10308
rect 11369 10364 11433 10368
rect 11369 10308 11373 10364
rect 11373 10308 11429 10364
rect 11429 10308 11433 10364
rect 11369 10304 11433 10308
rect 15200 10364 15264 10368
rect 15200 10308 15204 10364
rect 15204 10308 15260 10364
rect 15260 10308 15264 10364
rect 15200 10304 15264 10308
rect 15280 10364 15344 10368
rect 15280 10308 15284 10364
rect 15284 10308 15340 10364
rect 15340 10308 15344 10364
rect 15280 10304 15344 10308
rect 15360 10364 15424 10368
rect 15360 10308 15364 10364
rect 15364 10308 15420 10364
rect 15420 10308 15424 10364
rect 15360 10304 15424 10308
rect 15440 10364 15504 10368
rect 15440 10308 15444 10364
rect 15444 10308 15500 10364
rect 15500 10308 15504 10364
rect 15440 10304 15504 10308
rect 3647 9820 3711 9824
rect 3647 9764 3651 9820
rect 3651 9764 3707 9820
rect 3707 9764 3711 9820
rect 3647 9760 3711 9764
rect 3727 9820 3791 9824
rect 3727 9764 3731 9820
rect 3731 9764 3787 9820
rect 3787 9764 3791 9820
rect 3727 9760 3791 9764
rect 3807 9820 3871 9824
rect 3807 9764 3811 9820
rect 3811 9764 3867 9820
rect 3867 9764 3871 9820
rect 3807 9760 3871 9764
rect 3887 9820 3951 9824
rect 3887 9764 3891 9820
rect 3891 9764 3947 9820
rect 3947 9764 3951 9820
rect 3887 9760 3951 9764
rect 7718 9820 7782 9824
rect 7718 9764 7722 9820
rect 7722 9764 7778 9820
rect 7778 9764 7782 9820
rect 7718 9760 7782 9764
rect 7798 9820 7862 9824
rect 7798 9764 7802 9820
rect 7802 9764 7858 9820
rect 7858 9764 7862 9820
rect 7798 9760 7862 9764
rect 7878 9820 7942 9824
rect 7878 9764 7882 9820
rect 7882 9764 7938 9820
rect 7938 9764 7942 9820
rect 7878 9760 7942 9764
rect 7958 9820 8022 9824
rect 7958 9764 7962 9820
rect 7962 9764 8018 9820
rect 8018 9764 8022 9820
rect 7958 9760 8022 9764
rect 11789 9820 11853 9824
rect 11789 9764 11793 9820
rect 11793 9764 11849 9820
rect 11849 9764 11853 9820
rect 11789 9760 11853 9764
rect 11869 9820 11933 9824
rect 11869 9764 11873 9820
rect 11873 9764 11929 9820
rect 11929 9764 11933 9820
rect 11869 9760 11933 9764
rect 11949 9820 12013 9824
rect 11949 9764 11953 9820
rect 11953 9764 12009 9820
rect 12009 9764 12013 9820
rect 11949 9760 12013 9764
rect 12029 9820 12093 9824
rect 12029 9764 12033 9820
rect 12033 9764 12089 9820
rect 12089 9764 12093 9820
rect 12029 9760 12093 9764
rect 15860 9820 15924 9824
rect 15860 9764 15864 9820
rect 15864 9764 15920 9820
rect 15920 9764 15924 9820
rect 15860 9760 15924 9764
rect 15940 9820 16004 9824
rect 15940 9764 15944 9820
rect 15944 9764 16000 9820
rect 16000 9764 16004 9820
rect 15940 9760 16004 9764
rect 16020 9820 16084 9824
rect 16020 9764 16024 9820
rect 16024 9764 16080 9820
rect 16080 9764 16084 9820
rect 16020 9760 16084 9764
rect 16100 9820 16164 9824
rect 16100 9764 16104 9820
rect 16104 9764 16160 9820
rect 16160 9764 16164 9820
rect 16100 9760 16164 9764
rect 2987 9276 3051 9280
rect 2987 9220 2991 9276
rect 2991 9220 3047 9276
rect 3047 9220 3051 9276
rect 2987 9216 3051 9220
rect 3067 9276 3131 9280
rect 3067 9220 3071 9276
rect 3071 9220 3127 9276
rect 3127 9220 3131 9276
rect 3067 9216 3131 9220
rect 3147 9276 3211 9280
rect 3147 9220 3151 9276
rect 3151 9220 3207 9276
rect 3207 9220 3211 9276
rect 3147 9216 3211 9220
rect 3227 9276 3291 9280
rect 3227 9220 3231 9276
rect 3231 9220 3287 9276
rect 3287 9220 3291 9276
rect 3227 9216 3291 9220
rect 7058 9276 7122 9280
rect 7058 9220 7062 9276
rect 7062 9220 7118 9276
rect 7118 9220 7122 9276
rect 7058 9216 7122 9220
rect 7138 9276 7202 9280
rect 7138 9220 7142 9276
rect 7142 9220 7198 9276
rect 7198 9220 7202 9276
rect 7138 9216 7202 9220
rect 7218 9276 7282 9280
rect 7218 9220 7222 9276
rect 7222 9220 7278 9276
rect 7278 9220 7282 9276
rect 7218 9216 7282 9220
rect 7298 9276 7362 9280
rect 7298 9220 7302 9276
rect 7302 9220 7358 9276
rect 7358 9220 7362 9276
rect 7298 9216 7362 9220
rect 11129 9276 11193 9280
rect 11129 9220 11133 9276
rect 11133 9220 11189 9276
rect 11189 9220 11193 9276
rect 11129 9216 11193 9220
rect 11209 9276 11273 9280
rect 11209 9220 11213 9276
rect 11213 9220 11269 9276
rect 11269 9220 11273 9276
rect 11209 9216 11273 9220
rect 11289 9276 11353 9280
rect 11289 9220 11293 9276
rect 11293 9220 11349 9276
rect 11349 9220 11353 9276
rect 11289 9216 11353 9220
rect 11369 9276 11433 9280
rect 11369 9220 11373 9276
rect 11373 9220 11429 9276
rect 11429 9220 11433 9276
rect 11369 9216 11433 9220
rect 15200 9276 15264 9280
rect 15200 9220 15204 9276
rect 15204 9220 15260 9276
rect 15260 9220 15264 9276
rect 15200 9216 15264 9220
rect 15280 9276 15344 9280
rect 15280 9220 15284 9276
rect 15284 9220 15340 9276
rect 15340 9220 15344 9276
rect 15280 9216 15344 9220
rect 15360 9276 15424 9280
rect 15360 9220 15364 9276
rect 15364 9220 15420 9276
rect 15420 9220 15424 9276
rect 15360 9216 15424 9220
rect 15440 9276 15504 9280
rect 15440 9220 15444 9276
rect 15444 9220 15500 9276
rect 15500 9220 15504 9276
rect 15440 9216 15504 9220
rect 3647 8732 3711 8736
rect 3647 8676 3651 8732
rect 3651 8676 3707 8732
rect 3707 8676 3711 8732
rect 3647 8672 3711 8676
rect 3727 8732 3791 8736
rect 3727 8676 3731 8732
rect 3731 8676 3787 8732
rect 3787 8676 3791 8732
rect 3727 8672 3791 8676
rect 3807 8732 3871 8736
rect 3807 8676 3811 8732
rect 3811 8676 3867 8732
rect 3867 8676 3871 8732
rect 3807 8672 3871 8676
rect 3887 8732 3951 8736
rect 3887 8676 3891 8732
rect 3891 8676 3947 8732
rect 3947 8676 3951 8732
rect 3887 8672 3951 8676
rect 7718 8732 7782 8736
rect 7718 8676 7722 8732
rect 7722 8676 7778 8732
rect 7778 8676 7782 8732
rect 7718 8672 7782 8676
rect 7798 8732 7862 8736
rect 7798 8676 7802 8732
rect 7802 8676 7858 8732
rect 7858 8676 7862 8732
rect 7798 8672 7862 8676
rect 7878 8732 7942 8736
rect 7878 8676 7882 8732
rect 7882 8676 7938 8732
rect 7938 8676 7942 8732
rect 7878 8672 7942 8676
rect 7958 8732 8022 8736
rect 7958 8676 7962 8732
rect 7962 8676 8018 8732
rect 8018 8676 8022 8732
rect 7958 8672 8022 8676
rect 11789 8732 11853 8736
rect 11789 8676 11793 8732
rect 11793 8676 11849 8732
rect 11849 8676 11853 8732
rect 11789 8672 11853 8676
rect 11869 8732 11933 8736
rect 11869 8676 11873 8732
rect 11873 8676 11929 8732
rect 11929 8676 11933 8732
rect 11869 8672 11933 8676
rect 11949 8732 12013 8736
rect 11949 8676 11953 8732
rect 11953 8676 12009 8732
rect 12009 8676 12013 8732
rect 11949 8672 12013 8676
rect 12029 8732 12093 8736
rect 12029 8676 12033 8732
rect 12033 8676 12089 8732
rect 12089 8676 12093 8732
rect 12029 8672 12093 8676
rect 15860 8732 15924 8736
rect 15860 8676 15864 8732
rect 15864 8676 15920 8732
rect 15920 8676 15924 8732
rect 15860 8672 15924 8676
rect 15940 8732 16004 8736
rect 15940 8676 15944 8732
rect 15944 8676 16000 8732
rect 16000 8676 16004 8732
rect 15940 8672 16004 8676
rect 16020 8732 16084 8736
rect 16020 8676 16024 8732
rect 16024 8676 16080 8732
rect 16080 8676 16084 8732
rect 16020 8672 16084 8676
rect 16100 8732 16164 8736
rect 16100 8676 16104 8732
rect 16104 8676 16160 8732
rect 16160 8676 16164 8732
rect 16100 8672 16164 8676
rect 2987 8188 3051 8192
rect 2987 8132 2991 8188
rect 2991 8132 3047 8188
rect 3047 8132 3051 8188
rect 2987 8128 3051 8132
rect 3067 8188 3131 8192
rect 3067 8132 3071 8188
rect 3071 8132 3127 8188
rect 3127 8132 3131 8188
rect 3067 8128 3131 8132
rect 3147 8188 3211 8192
rect 3147 8132 3151 8188
rect 3151 8132 3207 8188
rect 3207 8132 3211 8188
rect 3147 8128 3211 8132
rect 3227 8188 3291 8192
rect 3227 8132 3231 8188
rect 3231 8132 3287 8188
rect 3287 8132 3291 8188
rect 3227 8128 3291 8132
rect 7058 8188 7122 8192
rect 7058 8132 7062 8188
rect 7062 8132 7118 8188
rect 7118 8132 7122 8188
rect 7058 8128 7122 8132
rect 7138 8188 7202 8192
rect 7138 8132 7142 8188
rect 7142 8132 7198 8188
rect 7198 8132 7202 8188
rect 7138 8128 7202 8132
rect 7218 8188 7282 8192
rect 7218 8132 7222 8188
rect 7222 8132 7278 8188
rect 7278 8132 7282 8188
rect 7218 8128 7282 8132
rect 7298 8188 7362 8192
rect 7298 8132 7302 8188
rect 7302 8132 7358 8188
rect 7358 8132 7362 8188
rect 7298 8128 7362 8132
rect 11129 8188 11193 8192
rect 11129 8132 11133 8188
rect 11133 8132 11189 8188
rect 11189 8132 11193 8188
rect 11129 8128 11193 8132
rect 11209 8188 11273 8192
rect 11209 8132 11213 8188
rect 11213 8132 11269 8188
rect 11269 8132 11273 8188
rect 11209 8128 11273 8132
rect 11289 8188 11353 8192
rect 11289 8132 11293 8188
rect 11293 8132 11349 8188
rect 11349 8132 11353 8188
rect 11289 8128 11353 8132
rect 11369 8188 11433 8192
rect 11369 8132 11373 8188
rect 11373 8132 11429 8188
rect 11429 8132 11433 8188
rect 11369 8128 11433 8132
rect 15200 8188 15264 8192
rect 15200 8132 15204 8188
rect 15204 8132 15260 8188
rect 15260 8132 15264 8188
rect 15200 8128 15264 8132
rect 15280 8188 15344 8192
rect 15280 8132 15284 8188
rect 15284 8132 15340 8188
rect 15340 8132 15344 8188
rect 15280 8128 15344 8132
rect 15360 8188 15424 8192
rect 15360 8132 15364 8188
rect 15364 8132 15420 8188
rect 15420 8132 15424 8188
rect 15360 8128 15424 8132
rect 15440 8188 15504 8192
rect 15440 8132 15444 8188
rect 15444 8132 15500 8188
rect 15500 8132 15504 8188
rect 15440 8128 15504 8132
rect 3647 7644 3711 7648
rect 3647 7588 3651 7644
rect 3651 7588 3707 7644
rect 3707 7588 3711 7644
rect 3647 7584 3711 7588
rect 3727 7644 3791 7648
rect 3727 7588 3731 7644
rect 3731 7588 3787 7644
rect 3787 7588 3791 7644
rect 3727 7584 3791 7588
rect 3807 7644 3871 7648
rect 3807 7588 3811 7644
rect 3811 7588 3867 7644
rect 3867 7588 3871 7644
rect 3807 7584 3871 7588
rect 3887 7644 3951 7648
rect 3887 7588 3891 7644
rect 3891 7588 3947 7644
rect 3947 7588 3951 7644
rect 3887 7584 3951 7588
rect 7718 7644 7782 7648
rect 7718 7588 7722 7644
rect 7722 7588 7778 7644
rect 7778 7588 7782 7644
rect 7718 7584 7782 7588
rect 7798 7644 7862 7648
rect 7798 7588 7802 7644
rect 7802 7588 7858 7644
rect 7858 7588 7862 7644
rect 7798 7584 7862 7588
rect 7878 7644 7942 7648
rect 7878 7588 7882 7644
rect 7882 7588 7938 7644
rect 7938 7588 7942 7644
rect 7878 7584 7942 7588
rect 7958 7644 8022 7648
rect 7958 7588 7962 7644
rect 7962 7588 8018 7644
rect 8018 7588 8022 7644
rect 7958 7584 8022 7588
rect 11789 7644 11853 7648
rect 11789 7588 11793 7644
rect 11793 7588 11849 7644
rect 11849 7588 11853 7644
rect 11789 7584 11853 7588
rect 11869 7644 11933 7648
rect 11869 7588 11873 7644
rect 11873 7588 11929 7644
rect 11929 7588 11933 7644
rect 11869 7584 11933 7588
rect 11949 7644 12013 7648
rect 11949 7588 11953 7644
rect 11953 7588 12009 7644
rect 12009 7588 12013 7644
rect 11949 7584 12013 7588
rect 12029 7644 12093 7648
rect 12029 7588 12033 7644
rect 12033 7588 12089 7644
rect 12089 7588 12093 7644
rect 12029 7584 12093 7588
rect 15860 7644 15924 7648
rect 15860 7588 15864 7644
rect 15864 7588 15920 7644
rect 15920 7588 15924 7644
rect 15860 7584 15924 7588
rect 15940 7644 16004 7648
rect 15940 7588 15944 7644
rect 15944 7588 16000 7644
rect 16000 7588 16004 7644
rect 15940 7584 16004 7588
rect 16020 7644 16084 7648
rect 16020 7588 16024 7644
rect 16024 7588 16080 7644
rect 16080 7588 16084 7644
rect 16020 7584 16084 7588
rect 16100 7644 16164 7648
rect 16100 7588 16104 7644
rect 16104 7588 16160 7644
rect 16160 7588 16164 7644
rect 16100 7584 16164 7588
rect 2987 7100 3051 7104
rect 2987 7044 2991 7100
rect 2991 7044 3047 7100
rect 3047 7044 3051 7100
rect 2987 7040 3051 7044
rect 3067 7100 3131 7104
rect 3067 7044 3071 7100
rect 3071 7044 3127 7100
rect 3127 7044 3131 7100
rect 3067 7040 3131 7044
rect 3147 7100 3211 7104
rect 3147 7044 3151 7100
rect 3151 7044 3207 7100
rect 3207 7044 3211 7100
rect 3147 7040 3211 7044
rect 3227 7100 3291 7104
rect 3227 7044 3231 7100
rect 3231 7044 3287 7100
rect 3287 7044 3291 7100
rect 3227 7040 3291 7044
rect 7058 7100 7122 7104
rect 7058 7044 7062 7100
rect 7062 7044 7118 7100
rect 7118 7044 7122 7100
rect 7058 7040 7122 7044
rect 7138 7100 7202 7104
rect 7138 7044 7142 7100
rect 7142 7044 7198 7100
rect 7198 7044 7202 7100
rect 7138 7040 7202 7044
rect 7218 7100 7282 7104
rect 7218 7044 7222 7100
rect 7222 7044 7278 7100
rect 7278 7044 7282 7100
rect 7218 7040 7282 7044
rect 7298 7100 7362 7104
rect 7298 7044 7302 7100
rect 7302 7044 7358 7100
rect 7358 7044 7362 7100
rect 7298 7040 7362 7044
rect 11129 7100 11193 7104
rect 11129 7044 11133 7100
rect 11133 7044 11189 7100
rect 11189 7044 11193 7100
rect 11129 7040 11193 7044
rect 11209 7100 11273 7104
rect 11209 7044 11213 7100
rect 11213 7044 11269 7100
rect 11269 7044 11273 7100
rect 11209 7040 11273 7044
rect 11289 7100 11353 7104
rect 11289 7044 11293 7100
rect 11293 7044 11349 7100
rect 11349 7044 11353 7100
rect 11289 7040 11353 7044
rect 11369 7100 11433 7104
rect 11369 7044 11373 7100
rect 11373 7044 11429 7100
rect 11429 7044 11433 7100
rect 11369 7040 11433 7044
rect 15200 7100 15264 7104
rect 15200 7044 15204 7100
rect 15204 7044 15260 7100
rect 15260 7044 15264 7100
rect 15200 7040 15264 7044
rect 15280 7100 15344 7104
rect 15280 7044 15284 7100
rect 15284 7044 15340 7100
rect 15340 7044 15344 7100
rect 15280 7040 15344 7044
rect 15360 7100 15424 7104
rect 15360 7044 15364 7100
rect 15364 7044 15420 7100
rect 15420 7044 15424 7100
rect 15360 7040 15424 7044
rect 15440 7100 15504 7104
rect 15440 7044 15444 7100
rect 15444 7044 15500 7100
rect 15500 7044 15504 7100
rect 15440 7040 15504 7044
rect 3647 6556 3711 6560
rect 3647 6500 3651 6556
rect 3651 6500 3707 6556
rect 3707 6500 3711 6556
rect 3647 6496 3711 6500
rect 3727 6556 3791 6560
rect 3727 6500 3731 6556
rect 3731 6500 3787 6556
rect 3787 6500 3791 6556
rect 3727 6496 3791 6500
rect 3807 6556 3871 6560
rect 3807 6500 3811 6556
rect 3811 6500 3867 6556
rect 3867 6500 3871 6556
rect 3807 6496 3871 6500
rect 3887 6556 3951 6560
rect 3887 6500 3891 6556
rect 3891 6500 3947 6556
rect 3947 6500 3951 6556
rect 3887 6496 3951 6500
rect 7718 6556 7782 6560
rect 7718 6500 7722 6556
rect 7722 6500 7778 6556
rect 7778 6500 7782 6556
rect 7718 6496 7782 6500
rect 7798 6556 7862 6560
rect 7798 6500 7802 6556
rect 7802 6500 7858 6556
rect 7858 6500 7862 6556
rect 7798 6496 7862 6500
rect 7878 6556 7942 6560
rect 7878 6500 7882 6556
rect 7882 6500 7938 6556
rect 7938 6500 7942 6556
rect 7878 6496 7942 6500
rect 7958 6556 8022 6560
rect 7958 6500 7962 6556
rect 7962 6500 8018 6556
rect 8018 6500 8022 6556
rect 7958 6496 8022 6500
rect 11789 6556 11853 6560
rect 11789 6500 11793 6556
rect 11793 6500 11849 6556
rect 11849 6500 11853 6556
rect 11789 6496 11853 6500
rect 11869 6556 11933 6560
rect 11869 6500 11873 6556
rect 11873 6500 11929 6556
rect 11929 6500 11933 6556
rect 11869 6496 11933 6500
rect 11949 6556 12013 6560
rect 11949 6500 11953 6556
rect 11953 6500 12009 6556
rect 12009 6500 12013 6556
rect 11949 6496 12013 6500
rect 12029 6556 12093 6560
rect 12029 6500 12033 6556
rect 12033 6500 12089 6556
rect 12089 6500 12093 6556
rect 12029 6496 12093 6500
rect 15860 6556 15924 6560
rect 15860 6500 15864 6556
rect 15864 6500 15920 6556
rect 15920 6500 15924 6556
rect 15860 6496 15924 6500
rect 15940 6556 16004 6560
rect 15940 6500 15944 6556
rect 15944 6500 16000 6556
rect 16000 6500 16004 6556
rect 15940 6496 16004 6500
rect 16020 6556 16084 6560
rect 16020 6500 16024 6556
rect 16024 6500 16080 6556
rect 16080 6500 16084 6556
rect 16020 6496 16084 6500
rect 16100 6556 16164 6560
rect 16100 6500 16104 6556
rect 16104 6500 16160 6556
rect 16160 6500 16164 6556
rect 16100 6496 16164 6500
rect 2987 6012 3051 6016
rect 2987 5956 2991 6012
rect 2991 5956 3047 6012
rect 3047 5956 3051 6012
rect 2987 5952 3051 5956
rect 3067 6012 3131 6016
rect 3067 5956 3071 6012
rect 3071 5956 3127 6012
rect 3127 5956 3131 6012
rect 3067 5952 3131 5956
rect 3147 6012 3211 6016
rect 3147 5956 3151 6012
rect 3151 5956 3207 6012
rect 3207 5956 3211 6012
rect 3147 5952 3211 5956
rect 3227 6012 3291 6016
rect 3227 5956 3231 6012
rect 3231 5956 3287 6012
rect 3287 5956 3291 6012
rect 3227 5952 3291 5956
rect 7058 6012 7122 6016
rect 7058 5956 7062 6012
rect 7062 5956 7118 6012
rect 7118 5956 7122 6012
rect 7058 5952 7122 5956
rect 7138 6012 7202 6016
rect 7138 5956 7142 6012
rect 7142 5956 7198 6012
rect 7198 5956 7202 6012
rect 7138 5952 7202 5956
rect 7218 6012 7282 6016
rect 7218 5956 7222 6012
rect 7222 5956 7278 6012
rect 7278 5956 7282 6012
rect 7218 5952 7282 5956
rect 7298 6012 7362 6016
rect 7298 5956 7302 6012
rect 7302 5956 7358 6012
rect 7358 5956 7362 6012
rect 7298 5952 7362 5956
rect 11129 6012 11193 6016
rect 11129 5956 11133 6012
rect 11133 5956 11189 6012
rect 11189 5956 11193 6012
rect 11129 5952 11193 5956
rect 11209 6012 11273 6016
rect 11209 5956 11213 6012
rect 11213 5956 11269 6012
rect 11269 5956 11273 6012
rect 11209 5952 11273 5956
rect 11289 6012 11353 6016
rect 11289 5956 11293 6012
rect 11293 5956 11349 6012
rect 11349 5956 11353 6012
rect 11289 5952 11353 5956
rect 11369 6012 11433 6016
rect 11369 5956 11373 6012
rect 11373 5956 11429 6012
rect 11429 5956 11433 6012
rect 11369 5952 11433 5956
rect 15200 6012 15264 6016
rect 15200 5956 15204 6012
rect 15204 5956 15260 6012
rect 15260 5956 15264 6012
rect 15200 5952 15264 5956
rect 15280 6012 15344 6016
rect 15280 5956 15284 6012
rect 15284 5956 15340 6012
rect 15340 5956 15344 6012
rect 15280 5952 15344 5956
rect 15360 6012 15424 6016
rect 15360 5956 15364 6012
rect 15364 5956 15420 6012
rect 15420 5956 15424 6012
rect 15360 5952 15424 5956
rect 15440 6012 15504 6016
rect 15440 5956 15444 6012
rect 15444 5956 15500 6012
rect 15500 5956 15504 6012
rect 15440 5952 15504 5956
rect 3647 5468 3711 5472
rect 3647 5412 3651 5468
rect 3651 5412 3707 5468
rect 3707 5412 3711 5468
rect 3647 5408 3711 5412
rect 3727 5468 3791 5472
rect 3727 5412 3731 5468
rect 3731 5412 3787 5468
rect 3787 5412 3791 5468
rect 3727 5408 3791 5412
rect 3807 5468 3871 5472
rect 3807 5412 3811 5468
rect 3811 5412 3867 5468
rect 3867 5412 3871 5468
rect 3807 5408 3871 5412
rect 3887 5468 3951 5472
rect 3887 5412 3891 5468
rect 3891 5412 3947 5468
rect 3947 5412 3951 5468
rect 3887 5408 3951 5412
rect 7718 5468 7782 5472
rect 7718 5412 7722 5468
rect 7722 5412 7778 5468
rect 7778 5412 7782 5468
rect 7718 5408 7782 5412
rect 7798 5468 7862 5472
rect 7798 5412 7802 5468
rect 7802 5412 7858 5468
rect 7858 5412 7862 5468
rect 7798 5408 7862 5412
rect 7878 5468 7942 5472
rect 7878 5412 7882 5468
rect 7882 5412 7938 5468
rect 7938 5412 7942 5468
rect 7878 5408 7942 5412
rect 7958 5468 8022 5472
rect 7958 5412 7962 5468
rect 7962 5412 8018 5468
rect 8018 5412 8022 5468
rect 7958 5408 8022 5412
rect 11789 5468 11853 5472
rect 11789 5412 11793 5468
rect 11793 5412 11849 5468
rect 11849 5412 11853 5468
rect 11789 5408 11853 5412
rect 11869 5468 11933 5472
rect 11869 5412 11873 5468
rect 11873 5412 11929 5468
rect 11929 5412 11933 5468
rect 11869 5408 11933 5412
rect 11949 5468 12013 5472
rect 11949 5412 11953 5468
rect 11953 5412 12009 5468
rect 12009 5412 12013 5468
rect 11949 5408 12013 5412
rect 12029 5468 12093 5472
rect 12029 5412 12033 5468
rect 12033 5412 12089 5468
rect 12089 5412 12093 5468
rect 12029 5408 12093 5412
rect 15860 5468 15924 5472
rect 15860 5412 15864 5468
rect 15864 5412 15920 5468
rect 15920 5412 15924 5468
rect 15860 5408 15924 5412
rect 15940 5468 16004 5472
rect 15940 5412 15944 5468
rect 15944 5412 16000 5468
rect 16000 5412 16004 5468
rect 15940 5408 16004 5412
rect 16020 5468 16084 5472
rect 16020 5412 16024 5468
rect 16024 5412 16080 5468
rect 16080 5412 16084 5468
rect 16020 5408 16084 5412
rect 16100 5468 16164 5472
rect 16100 5412 16104 5468
rect 16104 5412 16160 5468
rect 16160 5412 16164 5468
rect 16100 5408 16164 5412
rect 2987 4924 3051 4928
rect 2987 4868 2991 4924
rect 2991 4868 3047 4924
rect 3047 4868 3051 4924
rect 2987 4864 3051 4868
rect 3067 4924 3131 4928
rect 3067 4868 3071 4924
rect 3071 4868 3127 4924
rect 3127 4868 3131 4924
rect 3067 4864 3131 4868
rect 3147 4924 3211 4928
rect 3147 4868 3151 4924
rect 3151 4868 3207 4924
rect 3207 4868 3211 4924
rect 3147 4864 3211 4868
rect 3227 4924 3291 4928
rect 3227 4868 3231 4924
rect 3231 4868 3287 4924
rect 3287 4868 3291 4924
rect 3227 4864 3291 4868
rect 7058 4924 7122 4928
rect 7058 4868 7062 4924
rect 7062 4868 7118 4924
rect 7118 4868 7122 4924
rect 7058 4864 7122 4868
rect 7138 4924 7202 4928
rect 7138 4868 7142 4924
rect 7142 4868 7198 4924
rect 7198 4868 7202 4924
rect 7138 4864 7202 4868
rect 7218 4924 7282 4928
rect 7218 4868 7222 4924
rect 7222 4868 7278 4924
rect 7278 4868 7282 4924
rect 7218 4864 7282 4868
rect 7298 4924 7362 4928
rect 7298 4868 7302 4924
rect 7302 4868 7358 4924
rect 7358 4868 7362 4924
rect 7298 4864 7362 4868
rect 11129 4924 11193 4928
rect 11129 4868 11133 4924
rect 11133 4868 11189 4924
rect 11189 4868 11193 4924
rect 11129 4864 11193 4868
rect 11209 4924 11273 4928
rect 11209 4868 11213 4924
rect 11213 4868 11269 4924
rect 11269 4868 11273 4924
rect 11209 4864 11273 4868
rect 11289 4924 11353 4928
rect 11289 4868 11293 4924
rect 11293 4868 11349 4924
rect 11349 4868 11353 4924
rect 11289 4864 11353 4868
rect 11369 4924 11433 4928
rect 11369 4868 11373 4924
rect 11373 4868 11429 4924
rect 11429 4868 11433 4924
rect 11369 4864 11433 4868
rect 15200 4924 15264 4928
rect 15200 4868 15204 4924
rect 15204 4868 15260 4924
rect 15260 4868 15264 4924
rect 15200 4864 15264 4868
rect 15280 4924 15344 4928
rect 15280 4868 15284 4924
rect 15284 4868 15340 4924
rect 15340 4868 15344 4924
rect 15280 4864 15344 4868
rect 15360 4924 15424 4928
rect 15360 4868 15364 4924
rect 15364 4868 15420 4924
rect 15420 4868 15424 4924
rect 15360 4864 15424 4868
rect 15440 4924 15504 4928
rect 15440 4868 15444 4924
rect 15444 4868 15500 4924
rect 15500 4868 15504 4924
rect 15440 4864 15504 4868
rect 3647 4380 3711 4384
rect 3647 4324 3651 4380
rect 3651 4324 3707 4380
rect 3707 4324 3711 4380
rect 3647 4320 3711 4324
rect 3727 4380 3791 4384
rect 3727 4324 3731 4380
rect 3731 4324 3787 4380
rect 3787 4324 3791 4380
rect 3727 4320 3791 4324
rect 3807 4380 3871 4384
rect 3807 4324 3811 4380
rect 3811 4324 3867 4380
rect 3867 4324 3871 4380
rect 3807 4320 3871 4324
rect 3887 4380 3951 4384
rect 3887 4324 3891 4380
rect 3891 4324 3947 4380
rect 3947 4324 3951 4380
rect 3887 4320 3951 4324
rect 7718 4380 7782 4384
rect 7718 4324 7722 4380
rect 7722 4324 7778 4380
rect 7778 4324 7782 4380
rect 7718 4320 7782 4324
rect 7798 4380 7862 4384
rect 7798 4324 7802 4380
rect 7802 4324 7858 4380
rect 7858 4324 7862 4380
rect 7798 4320 7862 4324
rect 7878 4380 7942 4384
rect 7878 4324 7882 4380
rect 7882 4324 7938 4380
rect 7938 4324 7942 4380
rect 7878 4320 7942 4324
rect 7958 4380 8022 4384
rect 7958 4324 7962 4380
rect 7962 4324 8018 4380
rect 8018 4324 8022 4380
rect 7958 4320 8022 4324
rect 11789 4380 11853 4384
rect 11789 4324 11793 4380
rect 11793 4324 11849 4380
rect 11849 4324 11853 4380
rect 11789 4320 11853 4324
rect 11869 4380 11933 4384
rect 11869 4324 11873 4380
rect 11873 4324 11929 4380
rect 11929 4324 11933 4380
rect 11869 4320 11933 4324
rect 11949 4380 12013 4384
rect 11949 4324 11953 4380
rect 11953 4324 12009 4380
rect 12009 4324 12013 4380
rect 11949 4320 12013 4324
rect 12029 4380 12093 4384
rect 12029 4324 12033 4380
rect 12033 4324 12089 4380
rect 12089 4324 12093 4380
rect 12029 4320 12093 4324
rect 15860 4380 15924 4384
rect 15860 4324 15864 4380
rect 15864 4324 15920 4380
rect 15920 4324 15924 4380
rect 15860 4320 15924 4324
rect 15940 4380 16004 4384
rect 15940 4324 15944 4380
rect 15944 4324 16000 4380
rect 16000 4324 16004 4380
rect 15940 4320 16004 4324
rect 16020 4380 16084 4384
rect 16020 4324 16024 4380
rect 16024 4324 16080 4380
rect 16080 4324 16084 4380
rect 16020 4320 16084 4324
rect 16100 4380 16164 4384
rect 16100 4324 16104 4380
rect 16104 4324 16160 4380
rect 16160 4324 16164 4380
rect 16100 4320 16164 4324
rect 2987 3836 3051 3840
rect 2987 3780 2991 3836
rect 2991 3780 3047 3836
rect 3047 3780 3051 3836
rect 2987 3776 3051 3780
rect 3067 3836 3131 3840
rect 3067 3780 3071 3836
rect 3071 3780 3127 3836
rect 3127 3780 3131 3836
rect 3067 3776 3131 3780
rect 3147 3836 3211 3840
rect 3147 3780 3151 3836
rect 3151 3780 3207 3836
rect 3207 3780 3211 3836
rect 3147 3776 3211 3780
rect 3227 3836 3291 3840
rect 3227 3780 3231 3836
rect 3231 3780 3287 3836
rect 3287 3780 3291 3836
rect 3227 3776 3291 3780
rect 7058 3836 7122 3840
rect 7058 3780 7062 3836
rect 7062 3780 7118 3836
rect 7118 3780 7122 3836
rect 7058 3776 7122 3780
rect 7138 3836 7202 3840
rect 7138 3780 7142 3836
rect 7142 3780 7198 3836
rect 7198 3780 7202 3836
rect 7138 3776 7202 3780
rect 7218 3836 7282 3840
rect 7218 3780 7222 3836
rect 7222 3780 7278 3836
rect 7278 3780 7282 3836
rect 7218 3776 7282 3780
rect 7298 3836 7362 3840
rect 7298 3780 7302 3836
rect 7302 3780 7358 3836
rect 7358 3780 7362 3836
rect 7298 3776 7362 3780
rect 11129 3836 11193 3840
rect 11129 3780 11133 3836
rect 11133 3780 11189 3836
rect 11189 3780 11193 3836
rect 11129 3776 11193 3780
rect 11209 3836 11273 3840
rect 11209 3780 11213 3836
rect 11213 3780 11269 3836
rect 11269 3780 11273 3836
rect 11209 3776 11273 3780
rect 11289 3836 11353 3840
rect 11289 3780 11293 3836
rect 11293 3780 11349 3836
rect 11349 3780 11353 3836
rect 11289 3776 11353 3780
rect 11369 3836 11433 3840
rect 11369 3780 11373 3836
rect 11373 3780 11429 3836
rect 11429 3780 11433 3836
rect 11369 3776 11433 3780
rect 15200 3836 15264 3840
rect 15200 3780 15204 3836
rect 15204 3780 15260 3836
rect 15260 3780 15264 3836
rect 15200 3776 15264 3780
rect 15280 3836 15344 3840
rect 15280 3780 15284 3836
rect 15284 3780 15340 3836
rect 15340 3780 15344 3836
rect 15280 3776 15344 3780
rect 15360 3836 15424 3840
rect 15360 3780 15364 3836
rect 15364 3780 15420 3836
rect 15420 3780 15424 3836
rect 15360 3776 15424 3780
rect 15440 3836 15504 3840
rect 15440 3780 15444 3836
rect 15444 3780 15500 3836
rect 15500 3780 15504 3836
rect 15440 3776 15504 3780
rect 3647 3292 3711 3296
rect 3647 3236 3651 3292
rect 3651 3236 3707 3292
rect 3707 3236 3711 3292
rect 3647 3232 3711 3236
rect 3727 3292 3791 3296
rect 3727 3236 3731 3292
rect 3731 3236 3787 3292
rect 3787 3236 3791 3292
rect 3727 3232 3791 3236
rect 3807 3292 3871 3296
rect 3807 3236 3811 3292
rect 3811 3236 3867 3292
rect 3867 3236 3871 3292
rect 3807 3232 3871 3236
rect 3887 3292 3951 3296
rect 3887 3236 3891 3292
rect 3891 3236 3947 3292
rect 3947 3236 3951 3292
rect 3887 3232 3951 3236
rect 7718 3292 7782 3296
rect 7718 3236 7722 3292
rect 7722 3236 7778 3292
rect 7778 3236 7782 3292
rect 7718 3232 7782 3236
rect 7798 3292 7862 3296
rect 7798 3236 7802 3292
rect 7802 3236 7858 3292
rect 7858 3236 7862 3292
rect 7798 3232 7862 3236
rect 7878 3292 7942 3296
rect 7878 3236 7882 3292
rect 7882 3236 7938 3292
rect 7938 3236 7942 3292
rect 7878 3232 7942 3236
rect 7958 3292 8022 3296
rect 7958 3236 7962 3292
rect 7962 3236 8018 3292
rect 8018 3236 8022 3292
rect 7958 3232 8022 3236
rect 11789 3292 11853 3296
rect 11789 3236 11793 3292
rect 11793 3236 11849 3292
rect 11849 3236 11853 3292
rect 11789 3232 11853 3236
rect 11869 3292 11933 3296
rect 11869 3236 11873 3292
rect 11873 3236 11929 3292
rect 11929 3236 11933 3292
rect 11869 3232 11933 3236
rect 11949 3292 12013 3296
rect 11949 3236 11953 3292
rect 11953 3236 12009 3292
rect 12009 3236 12013 3292
rect 11949 3232 12013 3236
rect 12029 3292 12093 3296
rect 12029 3236 12033 3292
rect 12033 3236 12089 3292
rect 12089 3236 12093 3292
rect 12029 3232 12093 3236
rect 15860 3292 15924 3296
rect 15860 3236 15864 3292
rect 15864 3236 15920 3292
rect 15920 3236 15924 3292
rect 15860 3232 15924 3236
rect 15940 3292 16004 3296
rect 15940 3236 15944 3292
rect 15944 3236 16000 3292
rect 16000 3236 16004 3292
rect 15940 3232 16004 3236
rect 16020 3292 16084 3296
rect 16020 3236 16024 3292
rect 16024 3236 16080 3292
rect 16080 3236 16084 3292
rect 16020 3232 16084 3236
rect 16100 3292 16164 3296
rect 16100 3236 16104 3292
rect 16104 3236 16160 3292
rect 16160 3236 16164 3292
rect 16100 3232 16164 3236
rect 2987 2748 3051 2752
rect 2987 2692 2991 2748
rect 2991 2692 3047 2748
rect 3047 2692 3051 2748
rect 2987 2688 3051 2692
rect 3067 2748 3131 2752
rect 3067 2692 3071 2748
rect 3071 2692 3127 2748
rect 3127 2692 3131 2748
rect 3067 2688 3131 2692
rect 3147 2748 3211 2752
rect 3147 2692 3151 2748
rect 3151 2692 3207 2748
rect 3207 2692 3211 2748
rect 3147 2688 3211 2692
rect 3227 2748 3291 2752
rect 3227 2692 3231 2748
rect 3231 2692 3287 2748
rect 3287 2692 3291 2748
rect 3227 2688 3291 2692
rect 7058 2748 7122 2752
rect 7058 2692 7062 2748
rect 7062 2692 7118 2748
rect 7118 2692 7122 2748
rect 7058 2688 7122 2692
rect 7138 2748 7202 2752
rect 7138 2692 7142 2748
rect 7142 2692 7198 2748
rect 7198 2692 7202 2748
rect 7138 2688 7202 2692
rect 7218 2748 7282 2752
rect 7218 2692 7222 2748
rect 7222 2692 7278 2748
rect 7278 2692 7282 2748
rect 7218 2688 7282 2692
rect 7298 2748 7362 2752
rect 7298 2692 7302 2748
rect 7302 2692 7358 2748
rect 7358 2692 7362 2748
rect 7298 2688 7362 2692
rect 11129 2748 11193 2752
rect 11129 2692 11133 2748
rect 11133 2692 11189 2748
rect 11189 2692 11193 2748
rect 11129 2688 11193 2692
rect 11209 2748 11273 2752
rect 11209 2692 11213 2748
rect 11213 2692 11269 2748
rect 11269 2692 11273 2748
rect 11209 2688 11273 2692
rect 11289 2748 11353 2752
rect 11289 2692 11293 2748
rect 11293 2692 11349 2748
rect 11349 2692 11353 2748
rect 11289 2688 11353 2692
rect 11369 2748 11433 2752
rect 11369 2692 11373 2748
rect 11373 2692 11429 2748
rect 11429 2692 11433 2748
rect 11369 2688 11433 2692
rect 15200 2748 15264 2752
rect 15200 2692 15204 2748
rect 15204 2692 15260 2748
rect 15260 2692 15264 2748
rect 15200 2688 15264 2692
rect 15280 2748 15344 2752
rect 15280 2692 15284 2748
rect 15284 2692 15340 2748
rect 15340 2692 15344 2748
rect 15280 2688 15344 2692
rect 15360 2748 15424 2752
rect 15360 2692 15364 2748
rect 15364 2692 15420 2748
rect 15420 2692 15424 2748
rect 15360 2688 15424 2692
rect 15440 2748 15504 2752
rect 15440 2692 15444 2748
rect 15444 2692 15500 2748
rect 15500 2692 15504 2748
rect 15440 2688 15504 2692
rect 3647 2204 3711 2208
rect 3647 2148 3651 2204
rect 3651 2148 3707 2204
rect 3707 2148 3711 2204
rect 3647 2144 3711 2148
rect 3727 2204 3791 2208
rect 3727 2148 3731 2204
rect 3731 2148 3787 2204
rect 3787 2148 3791 2204
rect 3727 2144 3791 2148
rect 3807 2204 3871 2208
rect 3807 2148 3811 2204
rect 3811 2148 3867 2204
rect 3867 2148 3871 2204
rect 3807 2144 3871 2148
rect 3887 2204 3951 2208
rect 3887 2148 3891 2204
rect 3891 2148 3947 2204
rect 3947 2148 3951 2204
rect 3887 2144 3951 2148
rect 7718 2204 7782 2208
rect 7718 2148 7722 2204
rect 7722 2148 7778 2204
rect 7778 2148 7782 2204
rect 7718 2144 7782 2148
rect 7798 2204 7862 2208
rect 7798 2148 7802 2204
rect 7802 2148 7858 2204
rect 7858 2148 7862 2204
rect 7798 2144 7862 2148
rect 7878 2204 7942 2208
rect 7878 2148 7882 2204
rect 7882 2148 7938 2204
rect 7938 2148 7942 2204
rect 7878 2144 7942 2148
rect 7958 2204 8022 2208
rect 7958 2148 7962 2204
rect 7962 2148 8018 2204
rect 8018 2148 8022 2204
rect 7958 2144 8022 2148
rect 11789 2204 11853 2208
rect 11789 2148 11793 2204
rect 11793 2148 11849 2204
rect 11849 2148 11853 2204
rect 11789 2144 11853 2148
rect 11869 2204 11933 2208
rect 11869 2148 11873 2204
rect 11873 2148 11929 2204
rect 11929 2148 11933 2204
rect 11869 2144 11933 2148
rect 11949 2204 12013 2208
rect 11949 2148 11953 2204
rect 11953 2148 12009 2204
rect 12009 2148 12013 2204
rect 11949 2144 12013 2148
rect 12029 2204 12093 2208
rect 12029 2148 12033 2204
rect 12033 2148 12089 2204
rect 12089 2148 12093 2204
rect 12029 2144 12093 2148
rect 15860 2204 15924 2208
rect 15860 2148 15864 2204
rect 15864 2148 15920 2204
rect 15920 2148 15924 2204
rect 15860 2144 15924 2148
rect 15940 2204 16004 2208
rect 15940 2148 15944 2204
rect 15944 2148 16000 2204
rect 16000 2148 16004 2204
rect 15940 2144 16004 2148
rect 16020 2204 16084 2208
rect 16020 2148 16024 2204
rect 16024 2148 16080 2204
rect 16080 2148 16084 2204
rect 16020 2144 16084 2148
rect 16100 2204 16164 2208
rect 16100 2148 16104 2204
rect 16104 2148 16160 2204
rect 16160 2148 16164 2204
rect 16100 2144 16164 2148
<< metal4 >>
rect 2979 17984 3299 18000
rect 2979 17920 2987 17984
rect 3051 17920 3067 17984
rect 3131 17920 3147 17984
rect 3211 17920 3227 17984
rect 3291 17920 3299 17984
rect 2979 16896 3299 17920
rect 2979 16832 2987 16896
rect 3051 16832 3067 16896
rect 3131 16832 3147 16896
rect 3211 16832 3227 16896
rect 3291 16832 3299 16896
rect 2979 16098 3299 16832
rect 2979 15862 3021 16098
rect 3257 15862 3299 16098
rect 2979 15808 3299 15862
rect 2979 15744 2987 15808
rect 3051 15744 3067 15808
rect 3131 15744 3147 15808
rect 3211 15744 3227 15808
rect 3291 15744 3299 15808
rect 2979 14720 3299 15744
rect 2979 14656 2987 14720
rect 3051 14656 3067 14720
rect 3131 14656 3147 14720
rect 3211 14656 3227 14720
rect 3291 14656 3299 14720
rect 2979 13632 3299 14656
rect 2979 13568 2987 13632
rect 3051 13568 3067 13632
rect 3131 13568 3147 13632
rect 3211 13568 3227 13632
rect 3291 13568 3299 13632
rect 2979 12544 3299 13568
rect 2979 12480 2987 12544
rect 3051 12480 3067 12544
rect 3131 12480 3147 12544
rect 3211 12480 3227 12544
rect 3291 12480 3299 12544
rect 2979 12154 3299 12480
rect 2979 11918 3021 12154
rect 3257 11918 3299 12154
rect 2979 11456 3299 11918
rect 2979 11392 2987 11456
rect 3051 11392 3067 11456
rect 3131 11392 3147 11456
rect 3211 11392 3227 11456
rect 3291 11392 3299 11456
rect 2979 10368 3299 11392
rect 2979 10304 2987 10368
rect 3051 10304 3067 10368
rect 3131 10304 3147 10368
rect 3211 10304 3227 10368
rect 3291 10304 3299 10368
rect 2979 9280 3299 10304
rect 2979 9216 2987 9280
rect 3051 9216 3067 9280
rect 3131 9216 3147 9280
rect 3211 9216 3227 9280
rect 3291 9216 3299 9280
rect 2979 8210 3299 9216
rect 2979 8192 3021 8210
rect 3257 8192 3299 8210
rect 2979 8128 2987 8192
rect 3291 8128 3299 8192
rect 2979 7974 3021 8128
rect 3257 7974 3299 8128
rect 2979 7104 3299 7974
rect 2979 7040 2987 7104
rect 3051 7040 3067 7104
rect 3131 7040 3147 7104
rect 3211 7040 3227 7104
rect 3291 7040 3299 7104
rect 2979 6016 3299 7040
rect 2979 5952 2987 6016
rect 3051 5952 3067 6016
rect 3131 5952 3147 6016
rect 3211 5952 3227 6016
rect 3291 5952 3299 6016
rect 2979 4928 3299 5952
rect 2979 4864 2987 4928
rect 3051 4864 3067 4928
rect 3131 4864 3147 4928
rect 3211 4864 3227 4928
rect 3291 4864 3299 4928
rect 2979 4266 3299 4864
rect 2979 4030 3021 4266
rect 3257 4030 3299 4266
rect 2979 3840 3299 4030
rect 2979 3776 2987 3840
rect 3051 3776 3067 3840
rect 3131 3776 3147 3840
rect 3211 3776 3227 3840
rect 3291 3776 3299 3840
rect 2979 2752 3299 3776
rect 2979 2688 2987 2752
rect 3051 2688 3067 2752
rect 3131 2688 3147 2752
rect 3211 2688 3227 2752
rect 3291 2688 3299 2752
rect 2979 2128 3299 2688
rect 3639 17440 3959 18000
rect 3639 17376 3647 17440
rect 3711 17376 3727 17440
rect 3791 17376 3807 17440
rect 3871 17376 3887 17440
rect 3951 17376 3959 17440
rect 3639 16758 3959 17376
rect 3639 16522 3681 16758
rect 3917 16522 3959 16758
rect 3639 16352 3959 16522
rect 3639 16288 3647 16352
rect 3711 16288 3727 16352
rect 3791 16288 3807 16352
rect 3871 16288 3887 16352
rect 3951 16288 3959 16352
rect 3639 15264 3959 16288
rect 3639 15200 3647 15264
rect 3711 15200 3727 15264
rect 3791 15200 3807 15264
rect 3871 15200 3887 15264
rect 3951 15200 3959 15264
rect 3639 14176 3959 15200
rect 3639 14112 3647 14176
rect 3711 14112 3727 14176
rect 3791 14112 3807 14176
rect 3871 14112 3887 14176
rect 3951 14112 3959 14176
rect 3639 13088 3959 14112
rect 3639 13024 3647 13088
rect 3711 13024 3727 13088
rect 3791 13024 3807 13088
rect 3871 13024 3887 13088
rect 3951 13024 3959 13088
rect 3639 12814 3959 13024
rect 3639 12578 3681 12814
rect 3917 12578 3959 12814
rect 3639 12000 3959 12578
rect 3639 11936 3647 12000
rect 3711 11936 3727 12000
rect 3791 11936 3807 12000
rect 3871 11936 3887 12000
rect 3951 11936 3959 12000
rect 3639 10912 3959 11936
rect 3639 10848 3647 10912
rect 3711 10848 3727 10912
rect 3791 10848 3807 10912
rect 3871 10848 3887 10912
rect 3951 10848 3959 10912
rect 3639 9824 3959 10848
rect 3639 9760 3647 9824
rect 3711 9760 3727 9824
rect 3791 9760 3807 9824
rect 3871 9760 3887 9824
rect 3951 9760 3959 9824
rect 3639 8870 3959 9760
rect 3639 8736 3681 8870
rect 3917 8736 3959 8870
rect 3639 8672 3647 8736
rect 3951 8672 3959 8736
rect 3639 8634 3681 8672
rect 3917 8634 3959 8672
rect 3639 7648 3959 8634
rect 3639 7584 3647 7648
rect 3711 7584 3727 7648
rect 3791 7584 3807 7648
rect 3871 7584 3887 7648
rect 3951 7584 3959 7648
rect 3639 6560 3959 7584
rect 3639 6496 3647 6560
rect 3711 6496 3727 6560
rect 3791 6496 3807 6560
rect 3871 6496 3887 6560
rect 3951 6496 3959 6560
rect 3639 5472 3959 6496
rect 3639 5408 3647 5472
rect 3711 5408 3727 5472
rect 3791 5408 3807 5472
rect 3871 5408 3887 5472
rect 3951 5408 3959 5472
rect 3639 4926 3959 5408
rect 3639 4690 3681 4926
rect 3917 4690 3959 4926
rect 3639 4384 3959 4690
rect 3639 4320 3647 4384
rect 3711 4320 3727 4384
rect 3791 4320 3807 4384
rect 3871 4320 3887 4384
rect 3951 4320 3959 4384
rect 3639 3296 3959 4320
rect 3639 3232 3647 3296
rect 3711 3232 3727 3296
rect 3791 3232 3807 3296
rect 3871 3232 3887 3296
rect 3951 3232 3959 3296
rect 3639 2208 3959 3232
rect 3639 2144 3647 2208
rect 3711 2144 3727 2208
rect 3791 2144 3807 2208
rect 3871 2144 3887 2208
rect 3951 2144 3959 2208
rect 3639 2128 3959 2144
rect 7050 17984 7370 18000
rect 7050 17920 7058 17984
rect 7122 17920 7138 17984
rect 7202 17920 7218 17984
rect 7282 17920 7298 17984
rect 7362 17920 7370 17984
rect 7050 16896 7370 17920
rect 7050 16832 7058 16896
rect 7122 16832 7138 16896
rect 7202 16832 7218 16896
rect 7282 16832 7298 16896
rect 7362 16832 7370 16896
rect 7050 16098 7370 16832
rect 7050 15862 7092 16098
rect 7328 15862 7370 16098
rect 7050 15808 7370 15862
rect 7050 15744 7058 15808
rect 7122 15744 7138 15808
rect 7202 15744 7218 15808
rect 7282 15744 7298 15808
rect 7362 15744 7370 15808
rect 7050 14720 7370 15744
rect 7050 14656 7058 14720
rect 7122 14656 7138 14720
rect 7202 14656 7218 14720
rect 7282 14656 7298 14720
rect 7362 14656 7370 14720
rect 7050 13632 7370 14656
rect 7050 13568 7058 13632
rect 7122 13568 7138 13632
rect 7202 13568 7218 13632
rect 7282 13568 7298 13632
rect 7362 13568 7370 13632
rect 7050 12544 7370 13568
rect 7050 12480 7058 12544
rect 7122 12480 7138 12544
rect 7202 12480 7218 12544
rect 7282 12480 7298 12544
rect 7362 12480 7370 12544
rect 7050 12154 7370 12480
rect 7050 11918 7092 12154
rect 7328 11918 7370 12154
rect 7050 11456 7370 11918
rect 7050 11392 7058 11456
rect 7122 11392 7138 11456
rect 7202 11392 7218 11456
rect 7282 11392 7298 11456
rect 7362 11392 7370 11456
rect 7050 10368 7370 11392
rect 7050 10304 7058 10368
rect 7122 10304 7138 10368
rect 7202 10304 7218 10368
rect 7282 10304 7298 10368
rect 7362 10304 7370 10368
rect 7050 9280 7370 10304
rect 7050 9216 7058 9280
rect 7122 9216 7138 9280
rect 7202 9216 7218 9280
rect 7282 9216 7298 9280
rect 7362 9216 7370 9280
rect 7050 8210 7370 9216
rect 7050 8192 7092 8210
rect 7328 8192 7370 8210
rect 7050 8128 7058 8192
rect 7362 8128 7370 8192
rect 7050 7974 7092 8128
rect 7328 7974 7370 8128
rect 7050 7104 7370 7974
rect 7050 7040 7058 7104
rect 7122 7040 7138 7104
rect 7202 7040 7218 7104
rect 7282 7040 7298 7104
rect 7362 7040 7370 7104
rect 7050 6016 7370 7040
rect 7050 5952 7058 6016
rect 7122 5952 7138 6016
rect 7202 5952 7218 6016
rect 7282 5952 7298 6016
rect 7362 5952 7370 6016
rect 7050 4928 7370 5952
rect 7050 4864 7058 4928
rect 7122 4864 7138 4928
rect 7202 4864 7218 4928
rect 7282 4864 7298 4928
rect 7362 4864 7370 4928
rect 7050 4266 7370 4864
rect 7050 4030 7092 4266
rect 7328 4030 7370 4266
rect 7050 3840 7370 4030
rect 7050 3776 7058 3840
rect 7122 3776 7138 3840
rect 7202 3776 7218 3840
rect 7282 3776 7298 3840
rect 7362 3776 7370 3840
rect 7050 2752 7370 3776
rect 7050 2688 7058 2752
rect 7122 2688 7138 2752
rect 7202 2688 7218 2752
rect 7282 2688 7298 2752
rect 7362 2688 7370 2752
rect 7050 2128 7370 2688
rect 7710 17440 8030 18000
rect 7710 17376 7718 17440
rect 7782 17376 7798 17440
rect 7862 17376 7878 17440
rect 7942 17376 7958 17440
rect 8022 17376 8030 17440
rect 7710 16758 8030 17376
rect 7710 16522 7752 16758
rect 7988 16522 8030 16758
rect 7710 16352 8030 16522
rect 7710 16288 7718 16352
rect 7782 16288 7798 16352
rect 7862 16288 7878 16352
rect 7942 16288 7958 16352
rect 8022 16288 8030 16352
rect 7710 15264 8030 16288
rect 7710 15200 7718 15264
rect 7782 15200 7798 15264
rect 7862 15200 7878 15264
rect 7942 15200 7958 15264
rect 8022 15200 8030 15264
rect 7710 14176 8030 15200
rect 7710 14112 7718 14176
rect 7782 14112 7798 14176
rect 7862 14112 7878 14176
rect 7942 14112 7958 14176
rect 8022 14112 8030 14176
rect 7710 13088 8030 14112
rect 7710 13024 7718 13088
rect 7782 13024 7798 13088
rect 7862 13024 7878 13088
rect 7942 13024 7958 13088
rect 8022 13024 8030 13088
rect 7710 12814 8030 13024
rect 7710 12578 7752 12814
rect 7988 12578 8030 12814
rect 7710 12000 8030 12578
rect 7710 11936 7718 12000
rect 7782 11936 7798 12000
rect 7862 11936 7878 12000
rect 7942 11936 7958 12000
rect 8022 11936 8030 12000
rect 7710 10912 8030 11936
rect 7710 10848 7718 10912
rect 7782 10848 7798 10912
rect 7862 10848 7878 10912
rect 7942 10848 7958 10912
rect 8022 10848 8030 10912
rect 7710 9824 8030 10848
rect 7710 9760 7718 9824
rect 7782 9760 7798 9824
rect 7862 9760 7878 9824
rect 7942 9760 7958 9824
rect 8022 9760 8030 9824
rect 7710 8870 8030 9760
rect 7710 8736 7752 8870
rect 7988 8736 8030 8870
rect 7710 8672 7718 8736
rect 8022 8672 8030 8736
rect 7710 8634 7752 8672
rect 7988 8634 8030 8672
rect 7710 7648 8030 8634
rect 7710 7584 7718 7648
rect 7782 7584 7798 7648
rect 7862 7584 7878 7648
rect 7942 7584 7958 7648
rect 8022 7584 8030 7648
rect 7710 6560 8030 7584
rect 7710 6496 7718 6560
rect 7782 6496 7798 6560
rect 7862 6496 7878 6560
rect 7942 6496 7958 6560
rect 8022 6496 8030 6560
rect 7710 5472 8030 6496
rect 7710 5408 7718 5472
rect 7782 5408 7798 5472
rect 7862 5408 7878 5472
rect 7942 5408 7958 5472
rect 8022 5408 8030 5472
rect 7710 4926 8030 5408
rect 7710 4690 7752 4926
rect 7988 4690 8030 4926
rect 7710 4384 8030 4690
rect 7710 4320 7718 4384
rect 7782 4320 7798 4384
rect 7862 4320 7878 4384
rect 7942 4320 7958 4384
rect 8022 4320 8030 4384
rect 7710 3296 8030 4320
rect 7710 3232 7718 3296
rect 7782 3232 7798 3296
rect 7862 3232 7878 3296
rect 7942 3232 7958 3296
rect 8022 3232 8030 3296
rect 7710 2208 8030 3232
rect 7710 2144 7718 2208
rect 7782 2144 7798 2208
rect 7862 2144 7878 2208
rect 7942 2144 7958 2208
rect 8022 2144 8030 2208
rect 7710 2128 8030 2144
rect 11121 17984 11441 18000
rect 11121 17920 11129 17984
rect 11193 17920 11209 17984
rect 11273 17920 11289 17984
rect 11353 17920 11369 17984
rect 11433 17920 11441 17984
rect 11121 16896 11441 17920
rect 11121 16832 11129 16896
rect 11193 16832 11209 16896
rect 11273 16832 11289 16896
rect 11353 16832 11369 16896
rect 11433 16832 11441 16896
rect 11121 16098 11441 16832
rect 11121 15862 11163 16098
rect 11399 15862 11441 16098
rect 11121 15808 11441 15862
rect 11121 15744 11129 15808
rect 11193 15744 11209 15808
rect 11273 15744 11289 15808
rect 11353 15744 11369 15808
rect 11433 15744 11441 15808
rect 11121 14720 11441 15744
rect 11121 14656 11129 14720
rect 11193 14656 11209 14720
rect 11273 14656 11289 14720
rect 11353 14656 11369 14720
rect 11433 14656 11441 14720
rect 11121 13632 11441 14656
rect 11121 13568 11129 13632
rect 11193 13568 11209 13632
rect 11273 13568 11289 13632
rect 11353 13568 11369 13632
rect 11433 13568 11441 13632
rect 11121 12544 11441 13568
rect 11121 12480 11129 12544
rect 11193 12480 11209 12544
rect 11273 12480 11289 12544
rect 11353 12480 11369 12544
rect 11433 12480 11441 12544
rect 11121 12154 11441 12480
rect 11121 11918 11163 12154
rect 11399 11918 11441 12154
rect 11121 11456 11441 11918
rect 11121 11392 11129 11456
rect 11193 11392 11209 11456
rect 11273 11392 11289 11456
rect 11353 11392 11369 11456
rect 11433 11392 11441 11456
rect 11121 10368 11441 11392
rect 11121 10304 11129 10368
rect 11193 10304 11209 10368
rect 11273 10304 11289 10368
rect 11353 10304 11369 10368
rect 11433 10304 11441 10368
rect 11121 9280 11441 10304
rect 11121 9216 11129 9280
rect 11193 9216 11209 9280
rect 11273 9216 11289 9280
rect 11353 9216 11369 9280
rect 11433 9216 11441 9280
rect 11121 8210 11441 9216
rect 11121 8192 11163 8210
rect 11399 8192 11441 8210
rect 11121 8128 11129 8192
rect 11433 8128 11441 8192
rect 11121 7974 11163 8128
rect 11399 7974 11441 8128
rect 11121 7104 11441 7974
rect 11121 7040 11129 7104
rect 11193 7040 11209 7104
rect 11273 7040 11289 7104
rect 11353 7040 11369 7104
rect 11433 7040 11441 7104
rect 11121 6016 11441 7040
rect 11121 5952 11129 6016
rect 11193 5952 11209 6016
rect 11273 5952 11289 6016
rect 11353 5952 11369 6016
rect 11433 5952 11441 6016
rect 11121 4928 11441 5952
rect 11121 4864 11129 4928
rect 11193 4864 11209 4928
rect 11273 4864 11289 4928
rect 11353 4864 11369 4928
rect 11433 4864 11441 4928
rect 11121 4266 11441 4864
rect 11121 4030 11163 4266
rect 11399 4030 11441 4266
rect 11121 3840 11441 4030
rect 11121 3776 11129 3840
rect 11193 3776 11209 3840
rect 11273 3776 11289 3840
rect 11353 3776 11369 3840
rect 11433 3776 11441 3840
rect 11121 2752 11441 3776
rect 11121 2688 11129 2752
rect 11193 2688 11209 2752
rect 11273 2688 11289 2752
rect 11353 2688 11369 2752
rect 11433 2688 11441 2752
rect 11121 2128 11441 2688
rect 11781 17440 12101 18000
rect 11781 17376 11789 17440
rect 11853 17376 11869 17440
rect 11933 17376 11949 17440
rect 12013 17376 12029 17440
rect 12093 17376 12101 17440
rect 11781 16758 12101 17376
rect 11781 16522 11823 16758
rect 12059 16522 12101 16758
rect 11781 16352 12101 16522
rect 11781 16288 11789 16352
rect 11853 16288 11869 16352
rect 11933 16288 11949 16352
rect 12013 16288 12029 16352
rect 12093 16288 12101 16352
rect 11781 15264 12101 16288
rect 11781 15200 11789 15264
rect 11853 15200 11869 15264
rect 11933 15200 11949 15264
rect 12013 15200 12029 15264
rect 12093 15200 12101 15264
rect 11781 14176 12101 15200
rect 11781 14112 11789 14176
rect 11853 14112 11869 14176
rect 11933 14112 11949 14176
rect 12013 14112 12029 14176
rect 12093 14112 12101 14176
rect 11781 13088 12101 14112
rect 11781 13024 11789 13088
rect 11853 13024 11869 13088
rect 11933 13024 11949 13088
rect 12013 13024 12029 13088
rect 12093 13024 12101 13088
rect 11781 12814 12101 13024
rect 11781 12578 11823 12814
rect 12059 12578 12101 12814
rect 11781 12000 12101 12578
rect 11781 11936 11789 12000
rect 11853 11936 11869 12000
rect 11933 11936 11949 12000
rect 12013 11936 12029 12000
rect 12093 11936 12101 12000
rect 11781 10912 12101 11936
rect 11781 10848 11789 10912
rect 11853 10848 11869 10912
rect 11933 10848 11949 10912
rect 12013 10848 12029 10912
rect 12093 10848 12101 10912
rect 11781 9824 12101 10848
rect 11781 9760 11789 9824
rect 11853 9760 11869 9824
rect 11933 9760 11949 9824
rect 12013 9760 12029 9824
rect 12093 9760 12101 9824
rect 11781 8870 12101 9760
rect 11781 8736 11823 8870
rect 12059 8736 12101 8870
rect 11781 8672 11789 8736
rect 12093 8672 12101 8736
rect 11781 8634 11823 8672
rect 12059 8634 12101 8672
rect 11781 7648 12101 8634
rect 11781 7584 11789 7648
rect 11853 7584 11869 7648
rect 11933 7584 11949 7648
rect 12013 7584 12029 7648
rect 12093 7584 12101 7648
rect 11781 6560 12101 7584
rect 11781 6496 11789 6560
rect 11853 6496 11869 6560
rect 11933 6496 11949 6560
rect 12013 6496 12029 6560
rect 12093 6496 12101 6560
rect 11781 5472 12101 6496
rect 11781 5408 11789 5472
rect 11853 5408 11869 5472
rect 11933 5408 11949 5472
rect 12013 5408 12029 5472
rect 12093 5408 12101 5472
rect 11781 4926 12101 5408
rect 11781 4690 11823 4926
rect 12059 4690 12101 4926
rect 11781 4384 12101 4690
rect 11781 4320 11789 4384
rect 11853 4320 11869 4384
rect 11933 4320 11949 4384
rect 12013 4320 12029 4384
rect 12093 4320 12101 4384
rect 11781 3296 12101 4320
rect 11781 3232 11789 3296
rect 11853 3232 11869 3296
rect 11933 3232 11949 3296
rect 12013 3232 12029 3296
rect 12093 3232 12101 3296
rect 11781 2208 12101 3232
rect 11781 2144 11789 2208
rect 11853 2144 11869 2208
rect 11933 2144 11949 2208
rect 12013 2144 12029 2208
rect 12093 2144 12101 2208
rect 11781 2128 12101 2144
rect 15192 17984 15512 18000
rect 15192 17920 15200 17984
rect 15264 17920 15280 17984
rect 15344 17920 15360 17984
rect 15424 17920 15440 17984
rect 15504 17920 15512 17984
rect 15192 16896 15512 17920
rect 15192 16832 15200 16896
rect 15264 16832 15280 16896
rect 15344 16832 15360 16896
rect 15424 16832 15440 16896
rect 15504 16832 15512 16896
rect 15192 16098 15512 16832
rect 15192 15862 15234 16098
rect 15470 15862 15512 16098
rect 15192 15808 15512 15862
rect 15192 15744 15200 15808
rect 15264 15744 15280 15808
rect 15344 15744 15360 15808
rect 15424 15744 15440 15808
rect 15504 15744 15512 15808
rect 15192 14720 15512 15744
rect 15192 14656 15200 14720
rect 15264 14656 15280 14720
rect 15344 14656 15360 14720
rect 15424 14656 15440 14720
rect 15504 14656 15512 14720
rect 15192 13632 15512 14656
rect 15192 13568 15200 13632
rect 15264 13568 15280 13632
rect 15344 13568 15360 13632
rect 15424 13568 15440 13632
rect 15504 13568 15512 13632
rect 15192 12544 15512 13568
rect 15192 12480 15200 12544
rect 15264 12480 15280 12544
rect 15344 12480 15360 12544
rect 15424 12480 15440 12544
rect 15504 12480 15512 12544
rect 15192 12154 15512 12480
rect 15192 11918 15234 12154
rect 15470 11918 15512 12154
rect 15192 11456 15512 11918
rect 15192 11392 15200 11456
rect 15264 11392 15280 11456
rect 15344 11392 15360 11456
rect 15424 11392 15440 11456
rect 15504 11392 15512 11456
rect 15192 10368 15512 11392
rect 15192 10304 15200 10368
rect 15264 10304 15280 10368
rect 15344 10304 15360 10368
rect 15424 10304 15440 10368
rect 15504 10304 15512 10368
rect 15192 9280 15512 10304
rect 15192 9216 15200 9280
rect 15264 9216 15280 9280
rect 15344 9216 15360 9280
rect 15424 9216 15440 9280
rect 15504 9216 15512 9280
rect 15192 8210 15512 9216
rect 15192 8192 15234 8210
rect 15470 8192 15512 8210
rect 15192 8128 15200 8192
rect 15504 8128 15512 8192
rect 15192 7974 15234 8128
rect 15470 7974 15512 8128
rect 15192 7104 15512 7974
rect 15192 7040 15200 7104
rect 15264 7040 15280 7104
rect 15344 7040 15360 7104
rect 15424 7040 15440 7104
rect 15504 7040 15512 7104
rect 15192 6016 15512 7040
rect 15192 5952 15200 6016
rect 15264 5952 15280 6016
rect 15344 5952 15360 6016
rect 15424 5952 15440 6016
rect 15504 5952 15512 6016
rect 15192 4928 15512 5952
rect 15192 4864 15200 4928
rect 15264 4864 15280 4928
rect 15344 4864 15360 4928
rect 15424 4864 15440 4928
rect 15504 4864 15512 4928
rect 15192 4266 15512 4864
rect 15192 4030 15234 4266
rect 15470 4030 15512 4266
rect 15192 3840 15512 4030
rect 15192 3776 15200 3840
rect 15264 3776 15280 3840
rect 15344 3776 15360 3840
rect 15424 3776 15440 3840
rect 15504 3776 15512 3840
rect 15192 2752 15512 3776
rect 15192 2688 15200 2752
rect 15264 2688 15280 2752
rect 15344 2688 15360 2752
rect 15424 2688 15440 2752
rect 15504 2688 15512 2752
rect 15192 2128 15512 2688
rect 15852 17440 16172 18000
rect 15852 17376 15860 17440
rect 15924 17376 15940 17440
rect 16004 17376 16020 17440
rect 16084 17376 16100 17440
rect 16164 17376 16172 17440
rect 15852 16758 16172 17376
rect 15852 16522 15894 16758
rect 16130 16522 16172 16758
rect 15852 16352 16172 16522
rect 15852 16288 15860 16352
rect 15924 16288 15940 16352
rect 16004 16288 16020 16352
rect 16084 16288 16100 16352
rect 16164 16288 16172 16352
rect 15852 15264 16172 16288
rect 15852 15200 15860 15264
rect 15924 15200 15940 15264
rect 16004 15200 16020 15264
rect 16084 15200 16100 15264
rect 16164 15200 16172 15264
rect 15852 14176 16172 15200
rect 15852 14112 15860 14176
rect 15924 14112 15940 14176
rect 16004 14112 16020 14176
rect 16084 14112 16100 14176
rect 16164 14112 16172 14176
rect 15852 13088 16172 14112
rect 15852 13024 15860 13088
rect 15924 13024 15940 13088
rect 16004 13024 16020 13088
rect 16084 13024 16100 13088
rect 16164 13024 16172 13088
rect 15852 12814 16172 13024
rect 15852 12578 15894 12814
rect 16130 12578 16172 12814
rect 15852 12000 16172 12578
rect 15852 11936 15860 12000
rect 15924 11936 15940 12000
rect 16004 11936 16020 12000
rect 16084 11936 16100 12000
rect 16164 11936 16172 12000
rect 15852 10912 16172 11936
rect 15852 10848 15860 10912
rect 15924 10848 15940 10912
rect 16004 10848 16020 10912
rect 16084 10848 16100 10912
rect 16164 10848 16172 10912
rect 15852 9824 16172 10848
rect 15852 9760 15860 9824
rect 15924 9760 15940 9824
rect 16004 9760 16020 9824
rect 16084 9760 16100 9824
rect 16164 9760 16172 9824
rect 15852 8870 16172 9760
rect 15852 8736 15894 8870
rect 16130 8736 16172 8870
rect 15852 8672 15860 8736
rect 16164 8672 16172 8736
rect 15852 8634 15894 8672
rect 16130 8634 16172 8672
rect 15852 7648 16172 8634
rect 15852 7584 15860 7648
rect 15924 7584 15940 7648
rect 16004 7584 16020 7648
rect 16084 7584 16100 7648
rect 16164 7584 16172 7648
rect 15852 6560 16172 7584
rect 15852 6496 15860 6560
rect 15924 6496 15940 6560
rect 16004 6496 16020 6560
rect 16084 6496 16100 6560
rect 16164 6496 16172 6560
rect 15852 5472 16172 6496
rect 15852 5408 15860 5472
rect 15924 5408 15940 5472
rect 16004 5408 16020 5472
rect 16084 5408 16100 5472
rect 16164 5408 16172 5472
rect 15852 4926 16172 5408
rect 15852 4690 15894 4926
rect 16130 4690 16172 4926
rect 15852 4384 16172 4690
rect 15852 4320 15860 4384
rect 15924 4320 15940 4384
rect 16004 4320 16020 4384
rect 16084 4320 16100 4384
rect 16164 4320 16172 4384
rect 15852 3296 16172 4320
rect 15852 3232 15860 3296
rect 15924 3232 15940 3296
rect 16004 3232 16020 3296
rect 16084 3232 16100 3296
rect 16164 3232 16172 3296
rect 15852 2208 16172 3232
rect 15852 2144 15860 2208
rect 15924 2144 15940 2208
rect 16004 2144 16020 2208
rect 16084 2144 16100 2208
rect 16164 2144 16172 2208
rect 15852 2128 16172 2144
<< via4 >>
rect 3021 15862 3257 16098
rect 3021 11918 3257 12154
rect 3021 8192 3257 8210
rect 3021 8128 3051 8192
rect 3051 8128 3067 8192
rect 3067 8128 3131 8192
rect 3131 8128 3147 8192
rect 3147 8128 3211 8192
rect 3211 8128 3227 8192
rect 3227 8128 3257 8192
rect 3021 7974 3257 8128
rect 3021 4030 3257 4266
rect 3681 16522 3917 16758
rect 3681 12578 3917 12814
rect 3681 8736 3917 8870
rect 3681 8672 3711 8736
rect 3711 8672 3727 8736
rect 3727 8672 3791 8736
rect 3791 8672 3807 8736
rect 3807 8672 3871 8736
rect 3871 8672 3887 8736
rect 3887 8672 3917 8736
rect 3681 8634 3917 8672
rect 3681 4690 3917 4926
rect 7092 15862 7328 16098
rect 7092 11918 7328 12154
rect 7092 8192 7328 8210
rect 7092 8128 7122 8192
rect 7122 8128 7138 8192
rect 7138 8128 7202 8192
rect 7202 8128 7218 8192
rect 7218 8128 7282 8192
rect 7282 8128 7298 8192
rect 7298 8128 7328 8192
rect 7092 7974 7328 8128
rect 7092 4030 7328 4266
rect 7752 16522 7988 16758
rect 7752 12578 7988 12814
rect 7752 8736 7988 8870
rect 7752 8672 7782 8736
rect 7782 8672 7798 8736
rect 7798 8672 7862 8736
rect 7862 8672 7878 8736
rect 7878 8672 7942 8736
rect 7942 8672 7958 8736
rect 7958 8672 7988 8736
rect 7752 8634 7988 8672
rect 7752 4690 7988 4926
rect 11163 15862 11399 16098
rect 11163 11918 11399 12154
rect 11163 8192 11399 8210
rect 11163 8128 11193 8192
rect 11193 8128 11209 8192
rect 11209 8128 11273 8192
rect 11273 8128 11289 8192
rect 11289 8128 11353 8192
rect 11353 8128 11369 8192
rect 11369 8128 11399 8192
rect 11163 7974 11399 8128
rect 11163 4030 11399 4266
rect 11823 16522 12059 16758
rect 11823 12578 12059 12814
rect 11823 8736 12059 8870
rect 11823 8672 11853 8736
rect 11853 8672 11869 8736
rect 11869 8672 11933 8736
rect 11933 8672 11949 8736
rect 11949 8672 12013 8736
rect 12013 8672 12029 8736
rect 12029 8672 12059 8736
rect 11823 8634 12059 8672
rect 11823 4690 12059 4926
rect 15234 15862 15470 16098
rect 15234 11918 15470 12154
rect 15234 8192 15470 8210
rect 15234 8128 15264 8192
rect 15264 8128 15280 8192
rect 15280 8128 15344 8192
rect 15344 8128 15360 8192
rect 15360 8128 15424 8192
rect 15424 8128 15440 8192
rect 15440 8128 15470 8192
rect 15234 7974 15470 8128
rect 15234 4030 15470 4266
rect 15894 16522 16130 16758
rect 15894 12578 16130 12814
rect 15894 8736 16130 8870
rect 15894 8672 15924 8736
rect 15924 8672 15940 8736
rect 15940 8672 16004 8736
rect 16004 8672 16020 8736
rect 16020 8672 16084 8736
rect 16084 8672 16100 8736
rect 16100 8672 16130 8736
rect 15894 8634 16130 8672
rect 15894 4690 16130 4926
<< metal5 >>
rect 1056 16758 17436 16800
rect 1056 16522 3681 16758
rect 3917 16522 7752 16758
rect 7988 16522 11823 16758
rect 12059 16522 15894 16758
rect 16130 16522 17436 16758
rect 1056 16480 17436 16522
rect 1056 16098 17436 16140
rect 1056 15862 3021 16098
rect 3257 15862 7092 16098
rect 7328 15862 11163 16098
rect 11399 15862 15234 16098
rect 15470 15862 17436 16098
rect 1056 15820 17436 15862
rect 1056 12814 17436 12856
rect 1056 12578 3681 12814
rect 3917 12578 7752 12814
rect 7988 12578 11823 12814
rect 12059 12578 15894 12814
rect 16130 12578 17436 12814
rect 1056 12536 17436 12578
rect 1056 12154 17436 12196
rect 1056 11918 3021 12154
rect 3257 11918 7092 12154
rect 7328 11918 11163 12154
rect 11399 11918 15234 12154
rect 15470 11918 17436 12154
rect 1056 11876 17436 11918
rect 1056 8870 17436 8912
rect 1056 8634 3681 8870
rect 3917 8634 7752 8870
rect 7988 8634 11823 8870
rect 12059 8634 15894 8870
rect 16130 8634 17436 8870
rect 1056 8592 17436 8634
rect 1056 8210 17436 8252
rect 1056 7974 3021 8210
rect 3257 7974 7092 8210
rect 7328 7974 11163 8210
rect 11399 7974 15234 8210
rect 15470 7974 17436 8210
rect 1056 7932 17436 7974
rect 1056 4926 17436 4968
rect 1056 4690 3681 4926
rect 3917 4690 7752 4926
rect 7988 4690 11823 4926
rect 12059 4690 15894 4926
rect 16130 4690 17436 4926
rect 1056 4648 17436 4690
rect 1056 4266 17436 4308
rect 1056 4030 3021 4266
rect 3257 4030 7092 4266
rect 7328 4030 11163 4266
rect 11399 4030 15234 4266
rect 15470 4030 17436 4266
rect 1056 3988 17436 4030
use sky130_fd_sc_hd__clkbuf_4  _102_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 8556 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _103_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 7820 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _104_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 8004 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _105_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 8004 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _106_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 8832 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _107_
timestamp 1704896540
transform 1 0 10764 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _108_
timestamp 1704896540
transform -1 0 10212 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _109_
timestamp 1704896540
transform 1 0 10488 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _110_
timestamp 1704896540
transform 1 0 10488 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _111_
timestamp 1704896540
transform 1 0 9660 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _112_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 8924 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _113_
timestamp 1704896540
transform 1 0 10212 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _114_
timestamp 1704896540
transform -1 0 8832 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _115_
timestamp 1704896540
transform -1 0 8832 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _116_
timestamp 1704896540
transform 1 0 16100 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _117_
timestamp 1704896540
transform -1 0 16560 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _118_
timestamp 1704896540
transform -1 0 16652 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _119_
timestamp 1704896540
transform 1 0 15732 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _120_
timestamp 1704896540
transform 1 0 12328 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _121_
timestamp 1704896540
transform 1 0 13248 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _122_
timestamp 1704896540
transform -1 0 12512 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _123_
timestamp 1704896540
transform -1 0 12144 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _124_
timestamp 1704896540
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _125_
timestamp 1704896540
transform 1 0 14076 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _126_
timestamp 1704896540
transform 1 0 13156 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _127_
timestamp 1704896540
transform 1 0 13340 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _128_
timestamp 1704896540
transform 1 0 15916 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _129_
timestamp 1704896540
transform 1 0 16468 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _130_
timestamp 1704896540
transform -1 0 15824 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _131_
timestamp 1704896540
transform -1 0 15180 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _132_
timestamp 1704896540
transform 1 0 13248 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _133_
timestamp 1704896540
transform -1 0 13156 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _134_
timestamp 1704896540
transform 1 0 12880 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _135_
timestamp 1704896540
transform 1 0 12512 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _136_
timestamp 1704896540
transform 1 0 15916 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _137_
timestamp 1704896540
transform 1 0 16468 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _138_
timestamp 1704896540
transform -1 0 16008 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _139_
timestamp 1704896540
transform 1 0 15456 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _140_
timestamp 1704896540
transform 1 0 16008 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _141_
timestamp 1704896540
transform 1 0 16652 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _142_
timestamp 1704896540
transform -1 0 15824 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _143_
timestamp 1704896540
transform -1 0 15548 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _144_
timestamp 1704896540
transform 1 0 6072 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _145_
timestamp 1704896540
transform 1 0 14076 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _146_
timestamp 1704896540
transform -1 0 14076 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _147_
timestamp 1704896540
transform -1 0 13800 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _148_
timestamp 1704896540
transform 1 0 14076 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _149_
timestamp 1704896540
transform 1 0 11500 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _150_
timestamp 1704896540
transform -1 0 11408 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _151_
timestamp 1704896540
transform -1 0 10856 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _152_
timestamp 1704896540
transform 1 0 10304 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _153_
timestamp 1704896540
transform 1 0 9844 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _154_
timestamp 1704896540
transform 1 0 7728 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _155_
timestamp 1704896540
transform -1 0 10672 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _156_
timestamp 1704896540
transform 1 0 10396 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _157_
timestamp 1704896540
transform 1 0 10764 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _158_
timestamp 1704896540
transform -1 0 14628 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _159_
timestamp 1704896540
transform -1 0 14996 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _160_
timestamp 1704896540
transform 1 0 14812 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _161_
timestamp 1704896540
transform 1 0 15180 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _162_
timestamp 1704896540
transform -1 0 13432 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _163_
timestamp 1704896540
transform 1 0 13432 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _164_
timestamp 1704896540
transform -1 0 13524 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _165_
timestamp 1704896540
transform 1 0 14076 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _166_
timestamp 1704896540
transform -1 0 6256 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _167_
timestamp 1704896540
transform 1 0 6348 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _168_
timestamp 1704896540
transform -1 0 6624 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _169_
timestamp 1704896540
transform -1 0 6072 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _170_
timestamp 1704896540
transform 1 0 6072 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _171_
timestamp 1704896540
transform 1 0 6624 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _172_
timestamp 1704896540
transform 1 0 4968 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _173_
timestamp 1704896540
transform 1 0 5244 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _174_
timestamp 1704896540
transform 1 0 10672 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _175_
timestamp 1704896540
transform 1 0 11224 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _176_
timestamp 1704896540
transform -1 0 10488 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _177_
timestamp 1704896540
transform -1 0 10396 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _178_
timestamp 1704896540
transform 1 0 8280 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _179_
timestamp 1704896540
transform -1 0 8648 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _180_
timestamp 1704896540
transform -1 0 7912 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _181_
timestamp 1704896540
transform -1 0 7728 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _182_
timestamp 1704896540
transform 1 0 12052 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _183_
timestamp 1704896540
transform -1 0 12328 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _184_
timestamp 1704896540
transform 1 0 11592 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _185_
timestamp 1704896540
transform 1 0 10948 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _186_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 3588 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _187_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 3496 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _188_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 2576 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _189_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 4048 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _190_
timestamp 1704896540
transform 1 0 5612 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _191_
timestamp 1704896540
transform 1 0 5704 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _192_
timestamp 1704896540
transform -1 0 5060 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _193_
timestamp 1704896540
transform -1 0 4416 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _194_
timestamp 1704896540
transform 1 0 7820 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _195_
timestamp 1704896540
transform 1 0 8464 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _196_
timestamp 1704896540
transform -1 0 8280 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _197_
timestamp 1704896540
transform 1 0 8372 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _198_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 5244 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _199_
timestamp 1704896540
transform -1 0 7084 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _200_
timestamp 1704896540
transform -1 0 3496 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _201_
timestamp 1704896540
transform -1 0 5980 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _202_
timestamp 1704896540
transform -1 0 3496 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _203_
timestamp 1704896540
transform -1 0 9568 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _204_
timestamp 1704896540
transform -1 0 8280 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _205_
timestamp 1704896540
transform -1 0 2760 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _206_
timestamp 1704896540
transform -1 0 2484 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _207_
timestamp 1704896540
transform -1 0 7820 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _208_
timestamp 1704896540
transform -1 0 10488 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _209_
timestamp 1704896540
transform -1 0 9660 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _210_
timestamp 1704896540
transform -1 0 16284 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _211_
timestamp 1704896540
transform -1 0 12236 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _212_
timestamp 1704896540
transform -1 0 14076 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _213_
timestamp 1704896540
transform -1 0 15364 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _214_
timestamp 1704896540
transform -1 0 12880 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _215_
timestamp 1704896540
transform -1 0 15916 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _216_
timestamp 1704896540
transform -1 0 16652 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _217_
timestamp 1704896540
transform -1 0 14076 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _218_
timestamp 1704896540
transform -1 0 10580 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _219_
timestamp 1704896540
transform -1 0 10304 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _220_
timestamp 1704896540
transform -1 0 14812 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _221_
timestamp 1704896540
transform -1 0 14076 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _222_
timestamp 1704896540
transform -1 0 6348 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _223_
timestamp 1704896540
transform -1 0 5980 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _224_
timestamp 1704896540
transform -1 0 10672 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _225_
timestamp 1704896540
transform -1 0 8188 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _226_
timestamp 1704896540
transform 1 0 11224 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _227_
timestamp 1704896540
transform -1 0 5336 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _228_
timestamp 1704896540
transform -1 0 8372 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _229_
timestamp 1704896540
transform 1 0 5428 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _230_
timestamp 1704896540
transform 1 0 4876 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _231_
timestamp 1704896540
transform 1 0 4876 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _232_
timestamp 1704896540
transform 1 0 5612 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _233_
timestamp 1704896540
transform -1 0 6164 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _234_
timestamp 1704896540
transform 1 0 5244 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _235_
timestamp 1704896540
transform 1 0 6716 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _236_
timestamp 1704896540
transform 1 0 7268 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _237_
timestamp 1704896540
transform -1 0 7728 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _238_
timestamp 1704896540
transform 1 0 7084 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _239_
timestamp 1704896540
transform -1 0 3588 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _240_
timestamp 1704896540
transform 1 0 7176 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _241_
timestamp 1704896540
transform -1 0 2760 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _242_
timestamp 1704896540
transform 1 0 3312 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _243_
timestamp 1704896540
transform 1 0 3772 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _244_
timestamp 1704896540
transform -1 0 5612 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _245_
timestamp 1704896540
transform -1 0 5336 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _246_
timestamp 1704896540
transform -1 0 5612 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _247_
timestamp 1704896540
transform -1 0 6992 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _248_
timestamp 1704896540
transform -1 0 3588 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _249_
timestamp 1704896540
transform -1 0 2760 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _250_
timestamp 1704896540
transform 1 0 3404 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _251_
timestamp 1704896540
transform 1 0 3772 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _252_
timestamp 1704896540
transform -1 0 9476 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _253_
timestamp 1704896540
transform 1 0 8924 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _254_
timestamp 1704896540
transform 1 0 9476 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _255_
timestamp 1704896540
transform 1 0 9384 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _256_
timestamp 1704896540
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _257_
timestamp 1704896540
transform 1 0 8280 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _258_
timestamp 1704896540
transform -1 0 9476 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _259_
timestamp 1704896540
transform 1 0 8556 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _260_
timestamp 1704896540
transform 1 0 2668 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _261_
timestamp 1704896540
transform 1 0 3220 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _262_
timestamp 1704896540
transform -1 0 3036 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _263_
timestamp 1704896540
transform 1 0 3220 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _264_
timestamp 1704896540
transform 1 0 2484 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _265_
timestamp 1704896540
transform 1 0 3220 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _266_
timestamp 1704896540
transform -1 0 3312 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _267_
timestamp 1704896540
transform 1 0 1932 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__dfrtp_1  _268_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 1380 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _269_
timestamp 1704896540
transform -1 0 4416 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _270_
timestamp 1704896540
transform 1 0 1564 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _271_
timestamp 1704896540
transform 1 0 4232 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _272_
timestamp 1704896540
transform 1 0 5060 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _273_
timestamp 1704896540
transform 1 0 7912 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _274_
timestamp 1704896540
transform 1 0 9200 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _275_
timestamp 1704896540
transform 1 0 11500 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _276_
timestamp 1704896540
transform 1 0 12144 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _277_
timestamp 1704896540
transform 1 0 14260 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _278_
timestamp 1704896540
transform 1 0 14536 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _279_
timestamp 1704896540
transform -1 0 17112 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _280_
timestamp 1704896540
transform 1 0 14076 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _281_
timestamp 1704896540
transform -1 0 14444 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _282_
timestamp 1704896540
transform 1 0 10856 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _283_
timestamp 1704896540
transform -1 0 10856 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _284_
timestamp 1704896540
transform 1 0 8188 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _285_
timestamp 1704896540
transform -1 0 8188 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _286_
timestamp 1704896540
transform 1 0 3772 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _287_
timestamp 1704896540
transform 1 0 5980 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _288_
timestamp 1704896540
transform 1 0 6348 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _289_
timestamp 1704896540
transform 1 0 4416 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _290_
timestamp 1704896540
transform 1 0 3772 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _291_
timestamp 1704896540
transform -1 0 4784 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _292_
timestamp 1704896540
transform 1 0 1380 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _293_
timestamp 1704896540
transform 1 0 2576 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _294_
timestamp 1704896540
transform 1 0 4508 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _295_
timestamp 1704896540
transform 1 0 1380 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _296_
timestamp 1704896540
transform 1 0 1380 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _297_
timestamp 1704896540
transform 1 0 3772 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _298_
timestamp 1704896540
transform 1 0 4416 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _299_
timestamp 1704896540
transform 1 0 5796 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _300_
timestamp 1704896540
transform 1 0 6716 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _301_
timestamp 1704896540
transform 1 0 9292 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _302_
timestamp 1704896540
transform 1 0 11500 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _303_
timestamp 1704896540
transform -1 0 13340 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _304_
timestamp 1704896540
transform 1 0 6992 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _305_
timestamp 1704896540
transform 1 0 9568 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _306_
timestamp 1704896540
transform 1 0 9292 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _307_
timestamp 1704896540
transform -1 0 5612 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _308_
timestamp 1704896540
transform 1 0 1380 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _309_
timestamp 1704896540
transform 1 0 4416 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _310_
timestamp 1704896540
transform 1 0 3404 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _311_
timestamp 1704896540
transform 1 0 6164 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _312_
timestamp 1704896540
transform 1 0 7176 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _313_
timestamp 1704896540
transform 1 0 6900 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _314_
timestamp 1704896540
transform 1 0 6624 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _315_
timestamp 1704896540
transform 1 0 9108 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _316_
timestamp 1704896540
transform 1 0 8924 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _317_
timestamp 1704896540
transform 1 0 11500 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _318_
timestamp 1704896540
transform 1 0 11500 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _319_
timestamp 1704896540
transform 1 0 14076 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _320_
timestamp 1704896540
transform 1 0 14720 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _321_
timestamp 1704896540
transform -1 0 15640 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _322_
timestamp 1704896540
transform 1 0 8924 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _323_
timestamp 1704896540
transform 1 0 11500 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _324_
timestamp 1704896540
transform 1 0 11408 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _325_
timestamp 1704896540
transform 1 0 13340 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _326_
timestamp 1704896540
transform 1 0 11500 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _327_
timestamp 1704896540
transform 1 0 14260 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _328_
timestamp 1704896540
transform 1 0 14996 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _329_
timestamp 1704896540
transform -1 0 16560 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _330_
timestamp 1704896540
transform 1 0 13340 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _331_
timestamp 1704896540
transform 1 0 15272 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_4  fanout36
timestamp 1704896540
transform -1 0 7452 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout37 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 10396 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout38
timestamp 1704896540
transform -1 0 6900 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout39
timestamp 1704896540
transform -1 0 8464 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout40
timestamp 1704896540
transform 1 0 12696 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout41
timestamp 1704896540
transform -1 0 15732 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout42
timestamp 1704896540
transform -1 0 16192 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout43
timestamp 1704896540
transform -1 0 17020 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout44
timestamp 1704896540
transform -1 0 15548 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout45
timestamp 1704896540
transform -1 0 1748 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout46 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 7636 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  fanout47
timestamp 1704896540
transform 1 0 1472 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout48 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 6256 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout49
timestamp 1704896540
transform -1 0 9568 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  fanout50
timestamp 1704896540
transform 1 0 13064 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  fanout51
timestamp 1704896540
transform -1 0 10212 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout52
timestamp 1704896540
transform 1 0 13064 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  fanout53
timestamp 1704896540
transform 1 0 1564 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 1704896540
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 1704896540
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_41 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4876 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_48 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 5520 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_57
timestamp 1704896540
transform 1 0 6348 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_65
timestamp 1704896540
transform 1 0 7084 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_69
timestamp 1704896540
transform 1 0 7452 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_77 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 8188 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_83
timestamp 1704896540
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_85
timestamp 1704896540
transform 1 0 8924 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_93
timestamp 1704896540
transform 1 0 9660 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_97
timestamp 1704896540
transform 1 0 10028 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_104
timestamp 1704896540
transform 1 0 10672 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_111
timestamp 1704896540
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_120
timestamp 1704896540
transform 1 0 12144 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_128
timestamp 1704896540
transform 1 0 12880 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_132
timestamp 1704896540
transform 1 0 13248 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_141
timestamp 1704896540
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_153
timestamp 1704896540
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_165
timestamp 1704896540
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_169
timestamp 1704896540
transform 1 0 16652 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_173
timestamp 1704896540
transform 1 0 17020 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1704896540
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1704896540
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_27
timestamp 1704896540
transform 1 0 3588 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_35 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4324 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1704896540
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_84
timestamp 1704896540
transform 1 0 8832 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_106 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 10856 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_124
timestamp 1704896540
transform 1 0 12512 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_145
timestamp 1704896540
transform 1 0 14444 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_159
timestamp 1704896540
transform 1 0 15732 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 1704896540
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_169
timestamp 1704896540
transform 1 0 16652 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1704896540
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1704896540
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1704896540
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_73
timestamp 1704896540
transform 1 0 7820 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_103
timestamp 1704896540
transform 1 0 10580 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_136
timestamp 1704896540
transform 1 0 13616 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1704896540
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1704896540
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1704896540
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_39
timestamp 1704896540
transform 1 0 4692 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_47
timestamp 1704896540
transform 1 0 5428 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1704896540
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1704896540
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_69
timestamp 1704896540
transform 1 0 7452 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_101
timestamp 1704896540
transform 1 0 10396 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_109
timestamp 1704896540
transform 1 0 11132 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_113
timestamp 1704896540
transform 1 0 11500 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_121
timestamp 1704896540
transform 1 0 12236 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_128
timestamp 1704896540
transform 1 0 12880 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_140
timestamp 1704896540
transform 1 0 13984 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_160
timestamp 1704896540
transform 1 0 15824 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_169
timestamp 1704896540
transform 1 0 16652 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_173
timestamp 1704896540
transform 1 0 17020 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1704896540
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1704896540
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1704896540
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1704896540
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_41
timestamp 1704896540
transform 1 0 4876 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_72
timestamp 1704896540
transform 1 0 7728 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1704896540
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 1704896540
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_109
timestamp 1704896540
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_121
timestamp 1704896540
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_133
timestamp 1704896540
transform 1 0 13340 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_138
timestamp 1704896540
transform 1 0 13800 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_148
timestamp 1704896540
transform 1 0 14720 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_3
timestamp 1704896540
transform 1 0 1380 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_28
timestamp 1704896540
transform 1 0 3680 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_54
timestamp 1704896540
transform 1 0 6072 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_72
timestamp 1704896540
transform 1 0 7728 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_94
timestamp 1704896540
transform 1 0 9752 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_107
timestamp 1704896540
transform 1 0 10948 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1704896540
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_141
timestamp 1704896540
transform 1 0 14076 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_163
timestamp 1704896540
transform 1 0 16100 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_167
timestamp 1704896540
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_169
timestamp 1704896540
transform 1 0 16652 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_173
timestamp 1704896540
transform 1 0 17020 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_6
timestamp 1704896540
transform 1 0 1656 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_26
timestamp 1704896540
transform 1 0 3496 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_36
timestamp 1704896540
transform 1 0 4416 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_48
timestamp 1704896540
transform 1 0 5520 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_60
timestamp 1704896540
transform 1 0 6624 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_71
timestamp 1704896540
transform 1 0 7636 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1704896540
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_89
timestamp 1704896540
transform 1 0 9292 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_106
timestamp 1704896540
transform 1 0 10856 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_118
timestamp 1704896540
transform 1 0 11960 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_147
timestamp 1704896540
transform 1 0 14628 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_155
timestamp 1704896540
transform 1 0 15364 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_163
timestamp 1704896540
transform 1 0 16100 0 1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1704896540
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_15
timestamp 1704896540
transform 1 0 2484 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1704896540
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 1704896540
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 1704896540
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1704896540
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1704896540
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_69
timestamp 1704896540
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_87
timestamp 1704896540
transform 1 0 9108 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_119
timestamp 1704896540
transform 1 0 12052 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_131
timestamp 1704896540
transform 1 0 13156 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_141
timestamp 1704896540
transform 1 0 14076 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_153
timestamp 1704896540
transform 1 0 15180 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_162
timestamp 1704896540
transform 1 0 16008 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_169
timestamp 1704896540
transform 1 0 16652 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_173
timestamp 1704896540
transform 1 0 17020 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_26
timestamp 1704896540
transform 1 0 3496 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_32
timestamp 1704896540
transform 1 0 4048 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_40
timestamp 1704896540
transform 1 0 4784 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_51
timestamp 1704896540
transform 1 0 5796 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_60
timestamp 1704896540
transform 1 0 6624 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_64
timestamp 1704896540
transform 1 0 6992 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_79
timestamp 1704896540
transform 1 0 8372 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 1704896540
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_85
timestamp 1704896540
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_97
timestamp 1704896540
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_109
timestamp 1704896540
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_121
timestamp 1704896540
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 1704896540
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_141
timestamp 1704896540
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_171
timestamp 1704896540
transform 1 0 16836 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_3
timestamp 1704896540
transform 1 0 1380 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_11
timestamp 1704896540
transform 1 0 2116 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_84
timestamp 1704896540
transform 1 0 8832 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_92
timestamp 1704896540
transform 1 0 9568 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_99
timestamp 1704896540
transform 1 0 10212 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 1704896540
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_145
timestamp 1704896540
transform 1 0 14444 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_166
timestamp 1704896540
transform 1 0 16376 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_169
timestamp 1704896540
transform 1 0 16652 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_6
timestamp 1704896540
transform 1 0 1656 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_18
timestamp 1704896540
transform 1 0 2760 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1704896540
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1704896540
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 1704896540
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_53
timestamp 1704896540
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_65
timestamp 1704896540
transform 1 0 7084 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_78
timestamp 1704896540
transform 1 0 8280 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_111
timestamp 1704896540
transform 1 0 11316 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_123
timestamp 1704896540
transform 1 0 12420 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_134
timestamp 1704896540
transform 1 0 13432 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_141
timestamp 1704896540
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_153
timestamp 1704896540
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_165
timestamp 1704896540
transform 1 0 16284 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_9
timestamp 1704896540
transform 1 0 1932 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_17
timestamp 1704896540
transform 1 0 2668 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_40
timestamp 1704896540
transform 1 0 4784 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_46
timestamp 1704896540
transform 1 0 5336 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_54
timestamp 1704896540
transform 1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_61
timestamp 1704896540
transform 1 0 6716 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_79
timestamp 1704896540
transform 1 0 8372 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_91
timestamp 1704896540
transform 1 0 9476 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_105
timestamp 1704896540
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_111
timestamp 1704896540
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_140
timestamp 1704896540
transform 1 0 13984 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_169
timestamp 1704896540
transform 1 0 16652 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1704896540
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_85
timestamp 1704896540
transform 1 0 8924 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_92
timestamp 1704896540
transform 1 0 9568 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_100
timestamp 1704896540
transform 1 0 10304 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_109
timestamp 1704896540
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_121
timestamp 1704896540
transform 1 0 12236 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_129
timestamp 1704896540
transform 1 0 12972 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_173
timestamp 1704896540
transform 1 0 17020 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_24
timestamp 1704896540
transform 1 0 3312 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_36
timestamp 1704896540
transform 1 0 4416 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_48
timestamp 1704896540
transform 1 0 5520 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_57
timestamp 1704896540
transform 1 0 6348 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_86
timestamp 1704896540
transform 1 0 9016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_107
timestamp 1704896540
transform 1 0 10948 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_111
timestamp 1704896540
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_113
timestamp 1704896540
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_125
timestamp 1704896540
transform 1 0 12604 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_131
timestamp 1704896540
transform 1 0 13156 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_143
timestamp 1704896540
transform 1 0 14260 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_155
timestamp 1704896540
transform 1 0 15364 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_160
timestamp 1704896540
transform 1 0 15824 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_169
timestamp 1704896540
transform 1 0 16652 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_173
timestamp 1704896540
transform 1 0 17020 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_6
timestamp 1704896540
transform 1 0 1656 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_18
timestamp 1704896540
transform 1 0 2760 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_26
timestamp 1704896540
transform 1 0 3496 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_29
timestamp 1704896540
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_41
timestamp 1704896540
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_53
timestamp 1704896540
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_65
timestamp 1704896540
transform 1 0 7084 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_73
timestamp 1704896540
transform 1 0 7820 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_78
timestamp 1704896540
transform 1 0 8280 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_85
timestamp 1704896540
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_97
timestamp 1704896540
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_109
timestamp 1704896540
transform 1 0 11132 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_138
timestamp 1704896540
transform 1 0 13800 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_141
timestamp 1704896540
transform 1 0 14076 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_149
timestamp 1704896540
transform 1 0 14812 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_157
timestamp 1704896540
transform 1 0 15548 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_169
timestamp 1704896540
transform 1 0 16652 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_173
timestamp 1704896540
transform 1 0 17020 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_6
timestamp 1704896540
transform 1 0 1656 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_36
timestamp 1704896540
transform 1 0 4416 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_46
timestamp 1704896540
transform 1 0 5336 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_55
timestamp 1704896540
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_57
timestamp 1704896540
transform 1 0 6348 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_65
timestamp 1704896540
transform 1 0 7084 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_80
timestamp 1704896540
transform 1 0 8464 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_104
timestamp 1704896540
transform 1 0 10672 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_113
timestamp 1704896540
transform 1 0 11500 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_119
timestamp 1704896540
transform 1 0 12052 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_131
timestamp 1704896540
transform 1 0 13156 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_137
timestamp 1704896540
transform 1 0 13708 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_169
timestamp 1704896540
transform 1 0 16652 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_23
timestamp 1704896540
transform 1 0 3220 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 1704896540
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_36
timestamp 1704896540
transform 1 0 4416 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_83
timestamp 1704896540
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_112
timestamp 1704896540
transform 1 0 11408 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_131
timestamp 1704896540
transform 1 0 13156 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_139
timestamp 1704896540
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_141
timestamp 1704896540
transform 1 0 14076 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_149
timestamp 1704896540
transform 1 0 14812 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_3
timestamp 1704896540
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_15
timestamp 1704896540
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_27
timestamp 1704896540
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_39
timestamp 1704896540
transform 1 0 4692 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_43
timestamp 1704896540
transform 1 0 5060 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_49
timestamp 1704896540
transform 1 0 5612 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_54
timestamp 1704896540
transform 1 0 6072 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_57
timestamp 1704896540
transform 1 0 6348 0 -1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_72
timestamp 1704896540
transform 1 0 7728 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_84
timestamp 1704896540
transform 1 0 8832 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_92
timestamp 1704896540
transform 1 0 9568 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_104
timestamp 1704896540
transform 1 0 10672 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_153
timestamp 1704896540
transform 1 0 15180 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_173
timestamp 1704896540
transform 1 0 17020 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_3
timestamp 1704896540
transform 1 0 1380 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_9
timestamp 1704896540
transform 1 0 1932 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_21
timestamp 1704896540
transform 1 0 3036 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 1704896540
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_49
timestamp 1704896540
transform 1 0 5612 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_61
timestamp 1704896540
transform 1 0 6716 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_77
timestamp 1704896540
transform 1 0 8188 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_85
timestamp 1704896540
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_97
timestamp 1704896540
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_109
timestamp 1704896540
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_121
timestamp 1704896540
transform 1 0 12236 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_129
timestamp 1704896540
transform 1 0 12972 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_135
timestamp 1704896540
transform 1 0 13524 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_139
timestamp 1704896540
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_148
timestamp 1704896540
transform 1 0 14720 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_156
timestamp 1704896540
transform 1 0 15456 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_169
timestamp 1704896540
transform 1 0 16652 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_173
timestamp 1704896540
transform 1 0 17020 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_30
timestamp 1704896540
transform 1 0 3864 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_57
timestamp 1704896540
transform 1 0 6348 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_65
timestamp 1704896540
transform 1 0 7084 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_86
timestamp 1704896540
transform 1 0 9016 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_109
timestamp 1704896540
transform 1 0 11132 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_141
timestamp 1704896540
transform 1 0 14076 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_163
timestamp 1704896540
transform 1 0 16100 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_167
timestamp 1704896540
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_169
timestamp 1704896540
transform 1 0 16652 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_173
timestamp 1704896540
transform 1 0 17020 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_6
timestamp 1704896540
transform 1 0 1656 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_14
timestamp 1704896540
transform 1 0 2392 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 1704896540
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_29
timestamp 1704896540
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_41
timestamp 1704896540
transform 1 0 4876 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_53
timestamp 1704896540
transform 1 0 5980 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_64
timestamp 1704896540
transform 1 0 6992 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_70
timestamp 1704896540
transform 1 0 7544 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_74
timestamp 1704896540
transform 1 0 7912 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_82
timestamp 1704896540
transform 1 0 8648 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_85
timestamp 1704896540
transform 1 0 8924 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_93
timestamp 1704896540
transform 1 0 9660 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_114
timestamp 1704896540
transform 1 0 11592 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_126
timestamp 1704896540
transform 1 0 12696 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_138
timestamp 1704896540
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_141
timestamp 1704896540
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_153
timestamp 1704896540
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_165
timestamp 1704896540
transform 1 0 16284 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_6
timestamp 1704896540
transform 1 0 1656 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_18
timestamp 1704896540
transform 1 0 2760 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_30
timestamp 1704896540
transform 1 0 3864 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_42
timestamp 1704896540
transform 1 0 4968 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_52
timestamp 1704896540
transform 1 0 5888 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_57
timestamp 1704896540
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_69
timestamp 1704896540
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_81
timestamp 1704896540
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_93
timestamp 1704896540
transform 1 0 9660 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_102
timestamp 1704896540
transform 1 0 10488 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_110
timestamp 1704896540
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_113
timestamp 1704896540
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_125
timestamp 1704896540
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_137
timestamp 1704896540
transform 1 0 13708 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_145
timestamp 1704896540
transform 1 0 14444 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_169
timestamp 1704896540
transform 1 0 16652 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_3
timestamp 1704896540
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_15
timestamp 1704896540
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 1704896540
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_49
timestamp 1704896540
transform 1 0 5612 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_71
timestamp 1704896540
transform 1 0 7636 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_83
timestamp 1704896540
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_85
timestamp 1704896540
transform 1 0 8924 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_93
timestamp 1704896540
transform 1 0 9660 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_101
timestamp 1704896540
transform 1 0 10396 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_109
timestamp 1704896540
transform 1 0 11132 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_118
timestamp 1704896540
transform 1 0 11960 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_125
timestamp 1704896540
transform 1 0 12604 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_137
timestamp 1704896540
transform 1 0 13708 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_152
timestamp 1704896540
transform 1 0 15088 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_3
timestamp 1704896540
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_15
timestamp 1704896540
transform 1 0 2484 0 -1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_27
timestamp 1704896540
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_39
timestamp 1704896540
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_51
timestamp 1704896540
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_55
timestamp 1704896540
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_57
timestamp 1704896540
transform 1 0 6348 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_91
timestamp 1704896540
transform 1 0 9476 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_103
timestamp 1704896540
transform 1 0 10580 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_111
timestamp 1704896540
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_160
timestamp 1704896540
transform 1 0 15824 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_169
timestamp 1704896540
transform 1 0 16652 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_173
timestamp 1704896540
transform 1 0 17020 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_3
timestamp 1704896540
transform 1 0 1380 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_11
timestamp 1704896540
transform 1 0 2116 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_26
timestamp 1704896540
transform 1 0 3496 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_56
timestamp 1704896540
transform 1 0 6256 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_68
timestamp 1704896540
transform 1 0 7360 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_82
timestamp 1704896540
transform 1 0 8648 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_85
timestamp 1704896540
transform 1 0 8924 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_109
timestamp 1704896540
transform 1 0 11132 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_113
timestamp 1704896540
transform 1 0 11500 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_117
timestamp 1704896540
transform 1 0 11868 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_122
timestamp 1704896540
transform 1 0 12328 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_133
timestamp 1704896540
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_139
timestamp 1704896540
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_151
timestamp 1704896540
transform 1 0 14996 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_163
timestamp 1704896540
transform 1 0 16100 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_169
timestamp 1704896540
transform 1 0 16652 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_23
timestamp 1704896540
transform 1 0 3220 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_27
timestamp 1704896540
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_39
timestamp 1704896540
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_51
timestamp 1704896540
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_55
timestamp 1704896540
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_57
timestamp 1704896540
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_69
timestamp 1704896540
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_81
timestamp 1704896540
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_93
timestamp 1704896540
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_105
timestamp 1704896540
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_111
timestamp 1704896540
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_113
timestamp 1704896540
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_125
timestamp 1704896540
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_137
timestamp 1704896540
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_149
timestamp 1704896540
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_161
timestamp 1704896540
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_167
timestamp 1704896540
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_169
timestamp 1704896540
transform 1 0 16652 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_173
timestamp 1704896540
transform 1 0 17020 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_3
timestamp 1704896540
transform 1 0 1380 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_9
timestamp 1704896540
transform 1 0 1932 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_21
timestamp 1704896540
transform 1 0 3036 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_27
timestamp 1704896540
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_29
timestamp 1704896540
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_41
timestamp 1704896540
transform 1 0 4876 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_49
timestamp 1704896540
transform 1 0 5612 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_75
timestamp 1704896540
transform 1 0 8004 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_83
timestamp 1704896540
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_89
timestamp 1704896540
transform 1 0 9292 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_97
timestamp 1704896540
transform 1 0 10028 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_105
timestamp 1704896540
transform 1 0 10764 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_114
timestamp 1704896540
transform 1 0 11592 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_126
timestamp 1704896540
transform 1 0 12696 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_138
timestamp 1704896540
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_141
timestamp 1704896540
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_153
timestamp 1704896540
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_165
timestamp 1704896540
transform 1 0 16284 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_173
timestamp 1704896540
transform 1 0 17020 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_6
timestamp 1704896540
transform 1 0 1656 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_18
timestamp 1704896540
transform 1 0 2760 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_24
timestamp 1704896540
transform 1 0 3312 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_133
timestamp 1704896540
transform 1 0 13340 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_145
timestamp 1704896540
transform 1 0 14444 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_157
timestamp 1704896540
transform 1 0 15548 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_165
timestamp 1704896540
transform 1 0 16284 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_169
timestamp 1704896540
transform 1 0 16652 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_173
timestamp 1704896540
transform 1 0 17020 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_3
timestamp 1704896540
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_15
timestamp 1704896540
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_27
timestamp 1704896540
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_29
timestamp 1704896540
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_41
timestamp 1704896540
transform 1 0 4876 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_52
timestamp 1704896540
transform 1 0 5888 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_57
timestamp 1704896540
transform 1 0 6348 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_69
timestamp 1704896540
transform 1 0 7452 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_77
timestamp 1704896540
transform 1 0 8188 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_94
timestamp 1704896540
transform 1 0 9752 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_102
timestamp 1704896540
transform 1 0 10488 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_111
timestamp 1704896540
transform 1 0 11316 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_113
timestamp 1704896540
transform 1 0 11500 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_121
timestamp 1704896540
transform 1 0 12236 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_125
timestamp 1704896540
transform 1 0 12604 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_137
timestamp 1704896540
transform 1 0 13708 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_141
timestamp 1704896540
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_153
timestamp 1704896540
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_165
timestamp 1704896540
transform 1 0 16284 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_169
timestamp 1704896540
transform 1 0 16652 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_173
timestamp 1704896540
transform 1 0 17020 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1704896540
transform 1 0 16836 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1704896540
transform 1 0 5612 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1704896540
transform -1 0 2116 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 1704896540
transform 1 0 11040 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1704896540
transform 1 0 10212 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1704896540
transform -1 0 12604 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1704896540
transform -1 0 8556 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input8
timestamp 1704896540
transform 1 0 1380 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1704896540
transform -1 0 1656 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input10
timestamp 1704896540
transform 1 0 1380 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1704896540
transform -1 0 1656 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1704896540
transform 1 0 16836 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input13
timestamp 1704896540
transform 1 0 1656 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input14
timestamp 1704896540
transform -1 0 8740 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1704896540
transform -1 0 5520 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1704896540
transform -1 0 10028 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1704896540
transform -1 0 13248 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1704896540
transform 1 0 16836 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1704896540
transform 1 0 16836 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1704896540
transform 1 0 16836 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1704896540
transform -1 0 11316 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1704896540
transform -1 0 7452 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1704896540
transform 1 0 16836 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1704896540
transform -1 0 1656 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1704896540
transform -1 0 1656 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input26
timestamp 1704896540
transform -1 0 17112 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input27
timestamp 1704896540
transform -1 0 16560 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1704896540
transform 1 0 16836 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1704896540
transform 1 0 16836 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input30
timestamp 1704896540
transform 1 0 10396 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input31
timestamp 1704896540
transform 1 0 1380 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input32
timestamp 1704896540
transform -1 0 8832 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1704896540
transform -1 0 1656 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1704896540
transform 1 0 16836 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output35
timestamp 1704896540
transform -1 0 17112 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_29
timestamp 1704896540
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1704896540
transform -1 0 17388 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_30
timestamp 1704896540
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1704896540
transform -1 0 17388 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_31
timestamp 1704896540
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1704896540
transform -1 0 17388 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_32
timestamp 1704896540
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1704896540
transform -1 0 17388 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_33
timestamp 1704896540
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1704896540
transform -1 0 17388 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_34
timestamp 1704896540
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1704896540
transform -1 0 17388 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_35
timestamp 1704896540
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1704896540
transform -1 0 17388 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_36
timestamp 1704896540
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1704896540
transform -1 0 17388 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_37
timestamp 1704896540
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1704896540
transform -1 0 17388 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_38
timestamp 1704896540
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1704896540
transform -1 0 17388 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_39
timestamp 1704896540
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1704896540
transform -1 0 17388 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_40
timestamp 1704896540
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1704896540
transform -1 0 17388 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_41
timestamp 1704896540
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1704896540
transform -1 0 17388 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_42
timestamp 1704896540
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1704896540
transform -1 0 17388 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_43
timestamp 1704896540
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1704896540
transform -1 0 17388 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_44
timestamp 1704896540
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1704896540
transform -1 0 17388 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_45
timestamp 1704896540
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1704896540
transform -1 0 17388 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_46
timestamp 1704896540
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 1704896540
transform -1 0 17388 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_47
timestamp 1704896540
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 1704896540
transform -1 0 17388 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_48
timestamp 1704896540
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 1704896540
transform -1 0 17388 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_49
timestamp 1704896540
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 1704896540
transform -1 0 17388 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_50
timestamp 1704896540
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 1704896540
transform -1 0 17388 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_51
timestamp 1704896540
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 1704896540
transform -1 0 17388 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_52
timestamp 1704896540
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 1704896540
transform -1 0 17388 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_53
timestamp 1704896540
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 1704896540
transform -1 0 17388 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_54
timestamp 1704896540
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 1704896540
transform -1 0 17388 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_55
timestamp 1704896540
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 1704896540
transform -1 0 17388 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_56
timestamp 1704896540
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 1704896540
transform -1 0 17388 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_57
timestamp 1704896540
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp 1704896540
transform -1 0 17388 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_58 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_59
timestamp 1704896540
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_60
timestamp 1704896540
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_61
timestamp 1704896540
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_62
timestamp 1704896540
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_63
timestamp 1704896540
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_64
timestamp 1704896540
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_65
timestamp 1704896540
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_66
timestamp 1704896540
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_67
timestamp 1704896540
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_68
timestamp 1704896540
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_69
timestamp 1704896540
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_70
timestamp 1704896540
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_71
timestamp 1704896540
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_72
timestamp 1704896540
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_73
timestamp 1704896540
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_74
timestamp 1704896540
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_75
timestamp 1704896540
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_76
timestamp 1704896540
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_77
timestamp 1704896540
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_78
timestamp 1704896540
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_79
timestamp 1704896540
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_80
timestamp 1704896540
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_81
timestamp 1704896540
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_82
timestamp 1704896540
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_83
timestamp 1704896540
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_84
timestamp 1704896540
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_85
timestamp 1704896540
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_86
timestamp 1704896540
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_87
timestamp 1704896540
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_88
timestamp 1704896540
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_89
timestamp 1704896540
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_90
timestamp 1704896540
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_91
timestamp 1704896540
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_92
timestamp 1704896540
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_93
timestamp 1704896540
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_94
timestamp 1704896540
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_95
timestamp 1704896540
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_96
timestamp 1704896540
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_97
timestamp 1704896540
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_98
timestamp 1704896540
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_99
timestamp 1704896540
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_100
timestamp 1704896540
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_101
timestamp 1704896540
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_102
timestamp 1704896540
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_103
timestamp 1704896540
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_104
timestamp 1704896540
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_105
timestamp 1704896540
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_106
timestamp 1704896540
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_107
timestamp 1704896540
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_108
timestamp 1704896540
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_109
timestamp 1704896540
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_110
timestamp 1704896540
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_111
timestamp 1704896540
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_112
timestamp 1704896540
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_113
timestamp 1704896540
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_114
timestamp 1704896540
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_115
timestamp 1704896540
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_116
timestamp 1704896540
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_117
timestamp 1704896540
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_118
timestamp 1704896540
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_119
timestamp 1704896540
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_120
timestamp 1704896540
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_121
timestamp 1704896540
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_122
timestamp 1704896540
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_123
timestamp 1704896540
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_124
timestamp 1704896540
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_125
timestamp 1704896540
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_126
timestamp 1704896540
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_127
timestamp 1704896540
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_128
timestamp 1704896540
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_129
timestamp 1704896540
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_130
timestamp 1704896540
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_131
timestamp 1704896540
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_132
timestamp 1704896540
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_133
timestamp 1704896540
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_134
timestamp 1704896540
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_135
timestamp 1704896540
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_136
timestamp 1704896540
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_137
timestamp 1704896540
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_138
timestamp 1704896540
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_139
timestamp 1704896540
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_140
timestamp 1704896540
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_141
timestamp 1704896540
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_142
timestamp 1704896540
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_143
timestamp 1704896540
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_144
timestamp 1704896540
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_145
timestamp 1704896540
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_146
timestamp 1704896540
transform 1 0 6256 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_147
timestamp 1704896540
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_148
timestamp 1704896540
transform 1 0 11408 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_149
timestamp 1704896540
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_150
timestamp 1704896540
transform 1 0 16560 0 1 17408
box -38 -48 130 592
<< labels >>
flabel metal4 s 3639 2128 3959 18000 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 7710 2128 8030 18000 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 11781 2128 12101 18000 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 15852 2128 16172 18000 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 4648 17436 4968 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 8592 17436 8912 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 12536 17436 12856 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 16480 17436 16800 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 2979 2128 3299 18000 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 7050 2128 7370 18000 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 11121 2128 11441 18000 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 15192 2128 15512 18000 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 3988 17436 4308 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 7932 17436 8252 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 11876 17436 12196 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 15820 17436 16140 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 17716 14288 18516 14408 0 FreeSans 480 0 0 0 a[0]
port 2 nsew signal input
flabel metal2 s 5170 19860 5226 20660 0 FreeSans 224 90 0 0 a[10]
port 3 nsew signal input
flabel metal3 s 0 15648 800 15768 0 FreeSans 480 0 0 0 a[11]
port 4 nsew signal input
flabel metal2 s 10966 19860 11022 20660 0 FreeSans 224 90 0 0 a[12]
port 5 nsew signal input
flabel metal2 s 9678 19860 9734 20660 0 FreeSans 224 90 0 0 a[13]
port 6 nsew signal input
flabel metal2 s 12254 19860 12310 20660 0 FreeSans 224 90 0 0 a[14]
port 7 nsew signal input
flabel metal2 s 8390 19860 8446 20660 0 FreeSans 224 90 0 0 a[15]
port 8 nsew signal input
flabel metal3 s 0 12928 800 13048 0 FreeSans 480 0 0 0 a[16]
port 9 nsew signal input
flabel metal3 s 0 13608 800 13728 0 FreeSans 480 0 0 0 a[17]
port 10 nsew signal input
flabel metal3 s 0 10888 800 11008 0 FreeSans 480 0 0 0 a[18]
port 11 nsew signal input
flabel metal3 s 0 9528 800 9648 0 FreeSans 480 0 0 0 a[19]
port 12 nsew signal input
flabel metal3 s 17716 10888 18516 11008 0 FreeSans 480 0 0 0 a[1]
port 13 nsew signal input
flabel metal3 s 0 8168 800 8288 0 FreeSans 480 0 0 0 a[20]
port 14 nsew signal input
flabel metal2 s 8390 0 8446 800 0 FreeSans 224 90 0 0 a[21]
port 15 nsew signal input
flabel metal2 s 5170 0 5226 800 0 FreeSans 224 90 0 0 a[22]
port 16 nsew signal input
flabel metal2 s 9678 0 9734 800 0 FreeSans 224 90 0 0 a[23]
port 17 nsew signal input
flabel metal2 s 12898 0 12954 800 0 FreeSans 224 90 0 0 a[24]
port 18 nsew signal input
flabel metal3 s 17716 3408 18516 3528 0 FreeSans 480 0 0 0 a[25]
port 19 nsew signal input
flabel metal3 s 17716 6808 18516 6928 0 FreeSans 480 0 0 0 a[26]
port 20 nsew signal input
flabel metal3 s 17716 5448 18516 5568 0 FreeSans 480 0 0 0 a[27]
port 21 nsew signal input
flabel metal2 s 10966 0 11022 800 0 FreeSans 224 90 0 0 a[28]
port 22 nsew signal input
flabel metal2 s 7102 0 7158 800 0 FreeSans 224 90 0 0 a[29]
port 23 nsew signal input
flabel metal3 s 17716 12928 18516 13048 0 FreeSans 480 0 0 0 a[2]
port 24 nsew signal input
flabel metal3 s 0 5448 800 5568 0 FreeSans 480 0 0 0 a[30]
port 25 nsew signal input
flabel metal3 s 0 7488 800 7608 0 FreeSans 480 0 0 0 a[31]
port 26 nsew signal input
flabel metal3 s 17716 10208 18516 10328 0 FreeSans 480 0 0 0 a[3]
port 27 nsew signal input
flabel metal3 s 17716 11568 18516 11688 0 FreeSans 480 0 0 0 a[4]
port 28 nsew signal input
flabel metal3 s 17716 8848 18516 8968 0 FreeSans 480 0 0 0 a[5]
port 29 nsew signal input
flabel metal3 s 17716 7488 18516 7608 0 FreeSans 480 0 0 0 a[6]
port 30 nsew signal input
flabel metal2 s 10322 0 10378 800 0 FreeSans 224 90 0 0 a[7]
port 31 nsew signal input
flabel metal3 s 0 8848 800 8968 0 FreeSans 480 0 0 0 a[8]
port 32 nsew signal input
flabel metal2 s 9034 19860 9090 20660 0 FreeSans 224 90 0 0 a[9]
port 33 nsew signal input
flabel metal3 s 0 17008 800 17128 0 FreeSans 480 0 0 0 clk
port 34 nsew signal input
flabel metal3 s 17716 2728 18516 2848 0 FreeSans 480 0 0 0 rst
port 35 nsew signal input
flabel metal3 s 0 6808 800 6928 0 FreeSans 480 0 0 0 x
port 36 nsew signal input
flabel metal3 s 17716 14968 18516 15088 0 FreeSans 480 0 0 0 y
port 37 nsew signal output
rlabel metal1 9246 17408 9246 17408 0 VGND
rlabel metal1 9246 17952 9246 17952 0 VPWR
rlabel metal1 8464 6290 8464 6290 0 _000_
rlabel metal1 3220 13158 3220 13158 0 _001_
rlabel metal2 4738 3468 4738 3468 0 _002_
rlabel metal2 6118 3196 6118 3196 0 _003_
rlabel metal2 5382 2890 5382 2890 0 _004_
rlabel metal2 6578 4896 6578 4896 0 _005_
rlabel metal2 7038 5576 7038 5576 0 _006_
rlabel metal2 7590 4964 7590 4964 0 _007_
rlabel metal2 2990 15300 2990 15300 0 _008_
rlabel metal1 4554 17646 4554 17646 0 _009_
rlabel metal1 3036 15334 3036 15334 0 _010_
rlabel metal2 3910 15708 3910 15708 0 _011_
rlabel metal2 5474 17408 5474 17408 0 _012_
rlabel metal1 5566 17612 5566 17612 0 _013_
rlabel metal1 6670 17170 6670 17170 0 _014_
rlabel metal1 3174 5746 3174 5746 0 _015_
rlabel metal1 3450 5780 3450 5780 0 _016_
rlabel metal2 3542 5542 3542 5542 0 _017_
rlabel metal2 9430 17340 9430 17340 0 _018_
rlabel metal1 9384 17102 9384 17102 0 _019_
rlabel metal2 9522 17068 9522 17068 0 _020_
rlabel metal1 7912 14450 7912 14450 0 _021_
rlabel metal1 9016 15334 9016 15334 0 _022_
rlabel metal1 8878 14994 8878 14994 0 _023_
rlabel metal1 2622 12240 2622 12240 0 _024_
rlabel metal1 3220 12206 3220 12206 0 _025_
rlabel metal1 3128 12410 3128 12410 0 _026_
rlabel metal1 2714 9486 2714 9486 0 _027_
rlabel metal1 3312 9554 3312 9554 0 _028_
rlabel metal1 2254 10506 2254 10506 0 _029_
rlabel metal2 16330 5066 16330 5066 0 _030_
rlabel metal1 8050 6970 8050 6970 0 _031_
rlabel metal1 7636 7718 7636 7718 0 _032_
rlabel metal2 8510 7514 8510 7514 0 _033_
rlabel metal1 10718 8398 10718 8398 0 _034_
rlabel metal2 10442 7956 10442 7956 0 _035_
rlabel metal2 10626 8806 10626 8806 0 _036_
rlabel metal1 9430 3570 9430 3570 0 _037_
rlabel metal1 13570 3604 13570 3604 0 _038_
rlabel metal1 9706 3502 9706 3502 0 _039_
rlabel metal2 8694 3162 8694 3162 0 _040_
rlabel metal1 15686 11662 15686 11662 0 _041_
rlabel metal2 16238 11220 16238 11220 0 _042_
rlabel metal1 16192 12274 16192 12274 0 _043_
rlabel metal2 12282 3468 12282 3468 0 _044_
rlabel metal2 13386 3264 13386 3264 0 _045_
rlabel metal1 12190 2822 12190 2822 0 _046_
rlabel metal2 13570 7140 13570 7140 0 _047_
rlabel metal2 14030 7650 14030 7650 0 _048_
rlabel metal1 13386 8058 13386 8058 0 _049_
rlabel metal1 15870 3366 15870 3366 0 _050_
rlabel metal1 16192 4114 16192 4114 0 _051_
rlabel metal1 15364 4046 15364 4046 0 _052_
rlabel metal1 13110 10676 13110 10676 0 _053_
rlabel metal2 12834 10132 12834 10132 0 _054_
rlabel metal1 12926 10778 12926 10778 0 _055_
rlabel metal1 15410 6732 15410 6732 0 _056_
rlabel via1 16238 6834 16238 6834 0 _057_
rlabel metal2 15778 5916 15778 5916 0 _058_
rlabel metal1 15824 9486 15824 9486 0 _059_
rlabel metal1 16514 9010 16514 9010 0 _060_
rlabel metal1 15502 9690 15502 9690 0 _061_
rlabel metal1 11086 13328 11086 13328 0 _062_
rlabel metal1 13846 5202 13846 5202 0 _063_
rlabel metal2 14030 5712 14030 5712 0 _064_
rlabel metal1 13938 4658 13938 4658 0 _065_
rlabel metal2 10626 5882 10626 5882 0 _066_
rlabel metal2 10810 5916 10810 5916 0 _067_
rlabel metal2 10626 5338 10626 5338 0 _068_
rlabel metal1 9844 11526 9844 11526 0 _069_
rlabel metal1 12006 15538 12006 15538 0 _070_
rlabel metal2 10442 11254 10442 11254 0 _071_
rlabel metal2 10902 11356 10902 11356 0 _072_
rlabel metal1 14444 14450 14444 14450 0 _073_
rlabel metal2 14766 14892 14766 14892 0 _074_
rlabel metal2 14950 14756 14950 14756 0 _075_
rlabel metal2 13570 13056 13570 13056 0 _076_
rlabel metal1 13892 12954 13892 12954 0 _077_
rlabel metal1 13800 12342 13800 12342 0 _078_
rlabel metal2 6394 9146 6394 9146 0 _079_
rlabel metal2 6578 8772 6578 8772 0 _080_
rlabel metal1 6210 8398 6210 8398 0 _081_
rlabel metal1 5796 13362 5796 13362 0 _082_
rlabel metal1 6072 13294 6072 13294 0 _083_
rlabel metal1 5244 13498 5244 13498 0 _084_
rlabel metal1 10442 13294 10442 13294 0 _085_
rlabel metal1 10626 13396 10626 13396 0 _086_
rlabel metal2 10258 14246 10258 14246 0 _087_
rlabel metal1 7544 13294 7544 13294 0 _088_
rlabel metal1 7866 13328 7866 13328 0 _089_
rlabel metal1 7636 13158 7636 13158 0 _090_
rlabel metal2 11730 14960 11730 14960 0 _091_
rlabel metal1 11638 15436 11638 15436 0 _092_
rlabel metal1 11500 16626 11500 16626 0 _093_
rlabel metal1 3312 6766 3312 6766 0 _094_
rlabel metal1 3082 7208 3082 7208 0 _095_
rlabel metal1 4784 10574 4784 10574 0 _096_
rlabel metal1 5014 11696 5014 11696 0 _097_
rlabel metal2 4278 11356 4278 11356 0 _098_
rlabel metal1 8004 9554 8004 9554 0 _099_
rlabel metal2 8326 9316 8326 9316 0 _100_
rlabel metal2 8510 9690 8510 9690 0 _101_
rlabel metal2 17066 14127 17066 14127 0 a[0]
rlabel metal1 5842 17680 5842 17680 0 a[10]
rlabel metal3 866 15708 866 15708 0 a[11]
rlabel metal1 11040 17646 11040 17646 0 a[12]
rlabel metal1 10120 17646 10120 17646 0 a[13]
rlabel metal1 12328 17646 12328 17646 0 a[14]
rlabel metal1 8372 17646 8372 17646 0 a[15]
rlabel metal3 751 12988 751 12988 0 a[16]
rlabel metal3 1050 13668 1050 13668 0 a[17]
rlabel metal3 751 10948 751 10948 0 a[18]
rlabel metal3 1050 9588 1050 9588 0 a[19]
rlabel metal2 17066 11033 17066 11033 0 a[1]
rlabel metal3 1188 8228 1188 8228 0 a[20]
rlabel metal2 8418 1588 8418 1588 0 a[21]
rlabel metal2 5198 1588 5198 1588 0 a[22]
rlabel metal2 9706 1588 9706 1588 0 a[23]
rlabel metal2 12926 1588 12926 1588 0 a[24]
rlabel via2 17066 3485 17066 3485 0 a[25]
rlabel metal2 17066 7123 17066 7123 0 a[26]
rlabel metal2 17066 5593 17066 5593 0 a[27]
rlabel metal2 10994 1588 10994 1588 0 a[28]
rlabel metal2 7130 1588 7130 1588 0 a[29]
rlabel metal2 17066 13141 17066 13141 0 a[2]
rlabel metal3 1050 5508 1050 5508 0 a[30]
rlabel metal3 751 7548 751 7548 0 a[31]
rlabel metal2 17066 10455 17066 10455 0 a[3]
rlabel metal2 16514 11679 16514 11679 0 a[4]
rlabel metal2 17066 8687 17066 8687 0 a[5]
rlabel metal2 17066 7701 17066 7701 0 a[6]
rlabel metal2 10350 1588 10350 1588 0 a[7]
rlabel metal3 751 8908 751 8908 0 a[8]
rlabel metal1 8786 17680 8786 17680 0 a[9]
rlabel metal3 751 17068 751 17068 0 clk
rlabel metal1 2645 7378 2645 7378 0 dsa\[0\].last_carry
rlabel metal1 3634 6766 3634 6766 0 dsa\[0\].last_carry_next
rlabel metal1 2944 5678 2944 5678 0 dsa\[0\].y_out
rlabel metal1 4048 6970 4048 6970 0 dsa\[0\].y_out_next
rlabel metal2 8142 7650 8142 7650 0 dsa\[10\].last_carry
rlabel metal1 7038 6834 7038 6834 0 dsa\[10\].last_carry_next
rlabel metal1 7406 6698 7406 6698 0 dsa\[10\].y_in
rlabel metal1 6026 8466 6026 8466 0 dsa\[10\].y_out
rlabel metal1 8234 7208 8234 7208 0 dsa\[10\].y_out_next
rlabel metal2 5566 8670 5566 8670 0 dsa\[11\].last_carry
rlabel metal1 4876 9010 4876 9010 0 dsa\[11\].last_carry_next
rlabel metal2 2070 9044 2070 9044 0 dsa\[11\].y_out
rlabel metal1 5474 8432 5474 8432 0 dsa\[11\].y_out_next
rlabel metal2 2714 9350 2714 9350 0 dsa\[12\].last_carry
rlabel metal2 1702 9180 1702 9180 0 dsa\[12\].last_carry_next
rlabel metal1 4278 10778 4278 10778 0 dsa\[12\].y_out
rlabel metal1 2530 10744 2530 10744 0 dsa\[12\].y_out_next
rlabel metal1 6072 11322 6072 11322 0 dsa\[13\].last_carry
rlabel metal1 4738 10778 4738 10778 0 dsa\[13\].last_carry_next
rlabel metal1 2898 12784 2898 12784 0 dsa\[13\].y_out
rlabel metal1 2231 11186 2231 11186 0 dsa\[13\].y_out_next
rlabel metal2 3266 13090 3266 13090 0 dsa\[14\].last_carry
rlabel metal1 1886 12410 1886 12410 0 dsa\[14\].last_carry_next
rlabel metal1 5520 13906 5520 13906 0 dsa\[14\].y_out
rlabel metal1 3956 12682 3956 12682 0 dsa\[14\].y_out_next
rlabel metal2 6302 13124 6302 13124 0 dsa\[15\].last_carry
rlabel metal2 4738 13056 4738 13056 0 dsa\[15\].last_carry_next
rlabel metal1 7866 15436 7866 15436 0 dsa\[15\].y_out
rlabel metal1 5980 14042 5980 14042 0 dsa\[15\].y_out_next
rlabel metal1 8418 15130 8418 15130 0 dsa\[16\].last_carry
rlabel metal2 7038 15198 7038 15198 0 dsa\[16\].last_carry_next
rlabel metal1 11362 15334 11362 15334 0 dsa\[16\].y_out
rlabel metal1 9384 15130 9384 15130 0 dsa\[16\].y_out_next
rlabel metal2 12282 14892 12282 14892 0 dsa\[17\].last_carry
rlabel metal2 11914 14756 11914 14756 0 dsa\[17\].last_carry_next
rlabel metal1 9062 17102 9062 17102 0 dsa\[17\].y_out
rlabel metal2 13018 16932 13018 16932 0 dsa\[17\].y_out_next
rlabel via1 8970 17306 8970 17306 0 dsa\[18\].last_carry
rlabel metal1 8096 17102 8096 17102 0 dsa\[18\].last_carry_next
rlabel metal1 10856 16966 10856 16966 0 dsa\[18\].y_out
rlabel metal2 9890 16932 9890 16932 0 dsa\[18\].y_out_next
rlabel metal1 10902 13260 10902 13260 0 dsa\[19\].last_carry
rlabel metal2 9614 13022 9614 13022 0 dsa\[19\].last_carry_next
rlabel metal1 3542 15470 3542 15470 0 dsa\[19\].y_out
rlabel metal1 5290 14280 5290 14280 0 dsa\[19\].y_out_next
rlabel metal2 2898 5916 2898 5916 0 dsa\[1\].last_carry
rlabel metal1 1886 5304 1886 5304 0 dsa\[1\].last_carry_next
rlabel metal1 6670 5100 6670 5100 0 dsa\[1\].y_out
rlabel metal2 4554 5406 4554 5406 0 dsa\[1\].y_out_next
rlabel via1 2714 15419 2714 15419 0 dsa\[20\].last_carry
rlabel metal1 2254 15674 2254 15674 0 dsa\[20\].last_carry_next
rlabel metal2 6762 17119 6762 17119 0 dsa\[20\].y_out
rlabel metal1 4738 15368 4738 15368 0 dsa\[20\].y_out_next
rlabel metal1 5244 16966 5244 16966 0 dsa\[21\].last_carry
rlabel metal1 4508 17102 4508 17102 0 dsa\[21\].last_carry_next
rlabel metal2 8188 15164 8188 15164 0 dsa\[21\].y_out
rlabel metal2 6486 16796 6486 16796 0 dsa\[21\].y_out_next
rlabel metal2 8970 13090 8970 13090 0 dsa\[22\].last_carry
rlabel metal2 7498 12580 7498 12580 0 dsa\[22\].last_carry_next
rlabel metal1 8648 9554 8648 9554 0 dsa\[22\].y_out
rlabel metal1 7084 11186 7084 11186 0 dsa\[22\].y_out_next
rlabel metal2 8418 8670 8418 8670 0 dsa\[23\].last_carry
rlabel metal2 6946 9180 6946 9180 0 dsa\[23\].last_carry_next
rlabel metal2 10718 9146 10718 9146 0 dsa\[23\].y_out
rlabel metal1 9108 9418 9108 9418 0 dsa\[23\].y_out_next
rlabel metal2 10718 7582 10718 7582 0 dsa\[24\].last_carry
rlabel metal1 9522 7922 9522 7922 0 dsa\[24\].last_carry_next
rlabel metal1 13616 8466 13616 8466 0 dsa\[24\].y_out
rlabel metal1 11454 8534 11454 8534 0 dsa\[24\].y_out_next
rlabel metal1 13294 7480 13294 7480 0 dsa\[25\].last_carry
rlabel metal1 12604 7310 12604 7310 0 dsa\[25\].last_carry_next
rlabel metal1 15824 9146 15824 9146 0 dsa\[25\].y_out
rlabel metal2 13938 8738 13938 8738 0 dsa\[25\].y_out_next
rlabel metal1 16514 8942 16514 8942 0 dsa\[26\].last_carry
rlabel metal2 15042 8670 15042 8670 0 dsa\[26\].last_carry_next
rlabel metal2 10994 10812 10994 10812 0 dsa\[26\].y_out
rlabel metal1 14996 10234 14996 10234 0 dsa\[26\].y_out_next
rlabel metal2 10718 11492 10718 11492 0 dsa\[27\].last_carry
rlabel metal1 9430 10778 9430 10778 0 dsa\[27\].last_carry_next
rlabel metal1 13018 11118 13018 11118 0 dsa\[27\].y_out
rlabel metal1 11546 11322 11546 11322 0 dsa\[27\].y_out_next
rlabel metal1 13478 10064 13478 10064 0 dsa\[28\].last_carry
rlabel metal2 11730 10268 11730 10268 0 dsa\[28\].last_carry_next
rlabel metal1 13754 12750 13754 12750 0 dsa\[28\].y_out
rlabel metal1 13340 11322 13340 11322 0 dsa\[28\].y_out_next
rlabel metal2 13202 13124 13202 13124 0 dsa\[29\].last_carry
rlabel metal1 12604 12750 12604 12750 0 dsa\[29\].last_carry_next
rlabel metal1 16008 12206 16008 12206 0 dsa\[29\].y_out
rlabel metal2 14582 12580 14582 12580 0 dsa\[29\].y_out_next
rlabel metal2 6946 5236 6946 5236 0 dsa\[2\].last_carry
rlabel metal1 5888 4658 5888 4658 0 dsa\[2\].last_carry_next
rlabel metal2 10166 5508 10166 5508 0 dsa\[2\].y_out
rlabel metal1 7682 5304 7682 5304 0 dsa\[2\].y_out_next
rlabel metal2 16514 10948 16514 10948 0 dsa\[30\].last_carry
rlabel metal1 15502 11186 15502 11186 0 dsa\[30\].last_carry_next
rlabel metal2 14398 14654 14398 14654 0 dsa\[30\].y_out
rlabel via1 16244 13702 16244 13702 0 dsa\[30\].y_out_next
rlabel metal2 14950 15266 14950 15266 0 dsa\[31\].last_carry
rlabel metal2 14122 14756 14122 14756 0 dsa\[31\].last_carry_next
rlabel metal2 15594 14620 15594 14620 0 dsa\[31\].y_out_next
rlabel metal1 11362 6256 11362 6256 0 dsa\[3\].last_carry
rlabel metal2 9890 6052 9890 6052 0 dsa\[3\].last_carry_next
rlabel metal1 13662 5100 13662 5100 0 dsa\[3\].y_out
rlabel metal1 10902 5304 10902 5304 0 dsa\[3\].y_out_next
rlabel metal2 13938 6086 13938 6086 0 dsa\[4\].last_carry
rlabel metal1 12926 5338 12926 5338 0 dsa\[4\].last_carry_next
rlabel metal2 15686 6222 15686 6222 0 dsa\[4\].y_out
rlabel metal2 14582 4964 14582 4964 0 dsa\[4\].y_out_next
rlabel metal1 16238 6766 16238 6766 0 dsa\[5\].last_carry
rlabel metal1 15410 6834 15410 6834 0 dsa\[5\].last_carry_next
rlabel metal1 15134 4114 15134 4114 0 dsa\[5\].y_out
rlabel metal2 16790 5100 16790 5100 0 dsa\[5\].y_out_next
rlabel metal1 16146 3536 16146 3536 0 dsa\[6\].last_carry
rlabel metal2 14674 3298 14674 3298 0 dsa\[6\].last_carry_next
rlabel metal1 12535 2890 12535 2890 0 dsa\[6\].y_out
rlabel metal2 14122 3502 14122 3502 0 dsa\[6\].y_out_next
rlabel metal2 12650 3910 12650 3910 0 dsa\[7\].last_carry
rlabel metal1 11362 3162 11362 3162 0 dsa\[7\].last_carry_next
rlabel metal2 9062 3332 9062 3332 0 dsa\[7\].y_out
rlabel metal1 11132 2890 11132 2890 0 dsa\[7\].y_out_next
rlabel metal2 9890 3706 9890 3706 0 dsa\[8\].last_carry
rlabel metal2 8970 3876 8970 3876 0 dsa\[8\].last_carry_next
rlabel metal1 5474 2992 5474 2992 0 dsa\[8\].y_out
rlabel metal1 8234 3128 8234 3128 0 dsa\[8\].y_out_next
rlabel metal1 5336 3706 5336 3706 0 dsa\[9\].last_carry
rlabel metal1 4324 3162 4324 3162 0 dsa\[9\].last_carry_next
rlabel metal1 6072 3162 6072 3162 0 dsa\[9\].y_out_next
rlabel metal1 15686 15470 15686 15470 0 net1
rlabel metal1 2714 10540 2714 10540 0 net10
rlabel metal1 2300 9894 2300 9894 0 net11
rlabel metal1 16606 10642 16606 10642 0 net12
rlabel metal1 1886 8568 1886 8568 0 net13
rlabel metal1 8418 2618 8418 2618 0 net14
rlabel metal1 5566 3434 5566 3434 0 net15
rlabel metal1 10074 2618 10074 2618 0 net16
rlabel metal1 13340 2618 13340 2618 0 net17
rlabel metal1 16698 3400 16698 3400 0 net18
rlabel metal2 16698 6970 16698 6970 0 net19
rlabel metal1 5382 17782 5382 17782 0 net2
rlabel metal1 14582 5746 14582 5746 0 net20
rlabel metal1 11454 2618 11454 2618 0 net21
rlabel metal1 7130 5712 7130 5712 0 net22
rlabel metal1 15272 13226 15272 13226 0 net23
rlabel metal2 2530 5984 2530 5984 0 net24
rlabel metal2 2254 7718 2254 7718 0 net25
rlabel metal2 13754 10234 13754 10234 0 net26
rlabel metal1 15778 11866 15778 11866 0 net27
rlabel metal2 16882 9248 16882 9248 0 net28
rlabel metal2 14306 7582 14306 7582 0 net29
rlabel metal1 2300 15402 2300 15402 0 net3
rlabel metal1 10442 2618 10442 2618 0 net30
rlabel metal1 2185 8330 2185 8330 0 net31
rlabel metal1 8418 13328 8418 13328 0 net32
rlabel metal2 1610 16762 1610 16762 0 net33
rlabel metal1 16238 2890 16238 2890 0 net34
rlabel metal2 17066 15028 17066 15028 0 net35
rlabel metal1 6769 4522 6769 4522 0 net36
rlabel metal2 7314 7497 7314 7497 0 net37
rlabel metal1 3549 16150 3549 16150 0 net38
rlabel via1 8510 12869 8510 12869 0 net39
rlabel metal1 11408 17510 11408 17510 0 net4
rlabel metal2 12466 9248 12466 9248 0 net40
rlabel metal1 14805 3434 14805 3434 0 net41
rlabel metal1 10994 17129 10994 17129 0 net42
rlabel metal2 15686 14518 15686 14518 0 net43
rlabel metal1 16192 10710 16192 10710 0 net44
rlabel metal1 1610 5066 1610 5066 0 net45
rlabel metal1 6670 9078 6670 9078 0 net46
rlabel metal1 1610 15606 1610 15606 0 net47
rlabel metal1 6164 16626 6164 16626 0 net48
rlabel metal1 9200 9078 9200 9078 0 net49
rlabel metal2 8970 17714 8970 17714 0 net5
rlabel metal1 13754 8942 13754 8942 0 net50
rlabel metal1 11178 17850 11178 17850 0 net51
rlabel metal1 13340 14994 13340 14994 0 net52
rlabel metal1 6118 17170 6118 17170 0 net53
rlabel metal2 12558 16490 12558 16490 0 net6
rlabel metal1 8602 14382 8602 14382 0 net7
rlabel metal1 6486 13294 6486 13294 0 net8
rlabel metal1 3174 13328 3174 13328 0 net9
rlabel metal2 17066 2907 17066 2907 0 rst
rlabel metal2 4094 6817 4094 6817 0 x
rlabel metal2 16882 15181 16882 15181 0 y
<< properties >>
string FIXED_BBOX 0 0 18516 20660
<< end >>
