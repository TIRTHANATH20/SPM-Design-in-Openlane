VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO spm
  CLASS BLOCK ;
  FOREIGN spm ;
  ORIGIN 0.000 0.000 ;
  SIZE 92.580 BY 103.300 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 18.195 10.640 19.795 90.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 38.550 10.640 40.150 90.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 58.905 10.640 60.505 90.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 79.260 10.640 80.860 90.000 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 23.240 87.180 24.840 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 42.960 87.180 44.560 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 62.680 87.180 64.280 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 82.400 87.180 84.000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 14.895 10.640 16.495 90.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 35.250 10.640 36.850 90.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 55.605 10.640 57.205 90.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 75.960 10.640 77.560 90.000 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 19.940 87.180 21.540 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 39.660 87.180 41.260 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 59.380 87.180 60.980 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 79.100 87.180 80.700 ;
    END
  END VPWR
  PIN a[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 88.580 71.440 92.580 72.040 ;
    END
  END a[0]
  PIN a[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 25.850 99.300 26.130 103.300 ;
    END
  END a[10]
  PIN a[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 4.000 78.840 ;
    END
  END a[11]
  PIN a[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 54.830 99.300 55.110 103.300 ;
    END
  END a[12]
  PIN a[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 48.390 99.300 48.670 103.300 ;
    END
  END a[13]
  PIN a[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 61.270 99.300 61.550 103.300 ;
    END
  END a[14]
  PIN a[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 41.950 99.300 42.230 103.300 ;
    END
  END a[15]
  PIN a[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END a[16]
  PIN a[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END a[17]
  PIN a[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END a[18]
  PIN a[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END a[19]
  PIN a[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 88.580 54.440 92.580 55.040 ;
    END
  END a[1]
  PIN a[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END a[20]
  PIN a[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END a[21]
  PIN a[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END a[22]
  PIN a[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 4.000 ;
    END
  END a[23]
  PIN a[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END a[24]
  PIN a[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 88.580 17.040 92.580 17.640 ;
    END
  END a[25]
  PIN a[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 88.580 34.040 92.580 34.640 ;
    END
  END a[26]
  PIN a[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 88.580 27.240 92.580 27.840 ;
    END
  END a[27]
  PIN a[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 4.000 ;
    END
  END a[28]
  PIN a[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 4.000 ;
    END
  END a[29]
  PIN a[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 88.580 64.640 92.580 65.240 ;
    END
  END a[2]
  PIN a[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END a[30]
  PIN a[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END a[31]
  PIN a[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 88.580 51.040 92.580 51.640 ;
    END
  END a[3]
  PIN a[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 88.580 57.840 92.580 58.440 ;
    END
  END a[4]
  PIN a[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 88.580 44.240 92.580 44.840 ;
    END
  END a[5]
  PIN a[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 88.580 37.440 92.580 38.040 ;
    END
  END a[6]
  PIN a[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END a[7]
  PIN a[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END a[8]
  PIN a[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 45.170 99.300 45.450 103.300 ;
    END
  END a[9]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.040 4.000 85.640 ;
    END
  END clk
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 88.580 13.640 92.580 14.240 ;
    END
  END rst
  PIN x
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END x
  PIN y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 88.580 74.840 92.580 75.440 ;
    END
  END y
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 87.130 89.950 ;
      LAYER li1 ;
        RECT 5.520 10.795 86.940 89.845 ;
      LAYER met1 ;
        RECT 4.210 10.640 86.940 90.000 ;
      LAYER met2 ;
        RECT 4.230 99.020 25.570 99.300 ;
        RECT 26.410 99.020 41.670 99.300 ;
        RECT 42.510 99.020 44.890 99.300 ;
        RECT 45.730 99.020 48.110 99.300 ;
        RECT 48.950 99.020 54.550 99.300 ;
        RECT 55.390 99.020 60.990 99.300 ;
        RECT 61.830 99.020 85.470 99.300 ;
        RECT 4.230 4.280 85.470 99.020 ;
        RECT 4.230 4.000 25.570 4.280 ;
        RECT 26.410 4.000 35.230 4.280 ;
        RECT 36.070 4.000 41.670 4.280 ;
        RECT 42.510 4.000 48.110 4.280 ;
        RECT 48.950 4.000 51.330 4.280 ;
        RECT 52.170 4.000 54.550 4.280 ;
        RECT 55.390 4.000 64.210 4.280 ;
        RECT 65.050 4.000 85.470 4.280 ;
      LAYER met3 ;
        RECT 3.990 86.040 88.580 89.925 ;
        RECT 4.400 84.640 88.580 86.040 ;
        RECT 3.990 79.240 88.580 84.640 ;
        RECT 4.400 77.840 88.580 79.240 ;
        RECT 3.990 75.840 88.580 77.840 ;
        RECT 3.990 74.440 88.180 75.840 ;
        RECT 3.990 72.440 88.580 74.440 ;
        RECT 3.990 71.040 88.180 72.440 ;
        RECT 3.990 69.040 88.580 71.040 ;
        RECT 4.400 67.640 88.580 69.040 ;
        RECT 3.990 65.640 88.580 67.640 ;
        RECT 4.400 64.240 88.180 65.640 ;
        RECT 3.990 58.840 88.580 64.240 ;
        RECT 3.990 57.440 88.180 58.840 ;
        RECT 3.990 55.440 88.580 57.440 ;
        RECT 4.400 54.040 88.180 55.440 ;
        RECT 3.990 52.040 88.580 54.040 ;
        RECT 3.990 50.640 88.180 52.040 ;
        RECT 3.990 48.640 88.580 50.640 ;
        RECT 4.400 47.240 88.580 48.640 ;
        RECT 3.990 45.240 88.580 47.240 ;
        RECT 4.400 43.840 88.180 45.240 ;
        RECT 3.990 41.840 88.580 43.840 ;
        RECT 4.400 40.440 88.580 41.840 ;
        RECT 3.990 38.440 88.580 40.440 ;
        RECT 4.400 37.040 88.180 38.440 ;
        RECT 3.990 35.040 88.580 37.040 ;
        RECT 4.400 33.640 88.180 35.040 ;
        RECT 3.990 28.240 88.580 33.640 ;
        RECT 4.400 26.840 88.180 28.240 ;
        RECT 3.990 18.040 88.580 26.840 ;
        RECT 3.990 16.640 88.180 18.040 ;
        RECT 3.990 14.640 88.580 16.640 ;
        RECT 3.990 13.240 88.180 14.640 ;
        RECT 3.990 10.715 88.580 13.240 ;
  END
END spm
END LIBRARY

