magic
tech sky130A
magscale 1 2
timestamp 1742716875
<< nwell >>
rect 1066 2159 17426 17990
<< obsli1 >>
rect 1104 2159 17388 17969
<< obsm1 >>
rect 842 2128 17388 18000
<< metal2 >>
rect 5170 19860 5226 20660
rect 8390 19860 8446 20660
rect 9034 19860 9090 20660
rect 9678 19860 9734 20660
rect 10966 19860 11022 20660
rect 12254 19860 12310 20660
rect 5170 0 5226 800
rect 7102 0 7158 800
rect 8390 0 8446 800
rect 9678 0 9734 800
rect 10322 0 10378 800
rect 10966 0 11022 800
rect 12898 0 12954 800
<< obsm2 >>
rect 846 19804 5114 19860
rect 5282 19804 8334 19860
rect 8502 19804 8978 19860
rect 9146 19804 9622 19860
rect 9790 19804 10910 19860
rect 11078 19804 12198 19860
rect 12366 19804 17094 19860
rect 846 856 17094 19804
rect 846 800 5114 856
rect 5282 800 7046 856
rect 7214 800 8334 856
rect 8502 800 9622 856
rect 9790 800 10266 856
rect 10434 800 10910 856
rect 11078 800 12842 856
rect 13010 800 17094 856
<< metal3 >>
rect 0 17008 800 17128
rect 0 15648 800 15768
rect 17716 14968 18516 15088
rect 17716 14288 18516 14408
rect 0 13608 800 13728
rect 0 12928 800 13048
rect 17716 12928 18516 13048
rect 17716 11568 18516 11688
rect 0 10888 800 11008
rect 17716 10888 18516 11008
rect 17716 10208 18516 10328
rect 0 9528 800 9648
rect 0 8848 800 8968
rect 17716 8848 18516 8968
rect 0 8168 800 8288
rect 0 7488 800 7608
rect 17716 7488 18516 7608
rect 0 6808 800 6928
rect 17716 6808 18516 6928
rect 0 5448 800 5568
rect 17716 5448 18516 5568
rect 17716 3408 18516 3528
rect 17716 2728 18516 2848
<< obsm3 >>
rect 798 17208 17716 17985
rect 880 16928 17716 17208
rect 798 15848 17716 16928
rect 880 15568 17716 15848
rect 798 15168 17716 15568
rect 798 14888 17636 15168
rect 798 14488 17716 14888
rect 798 14208 17636 14488
rect 798 13808 17716 14208
rect 880 13528 17716 13808
rect 798 13128 17716 13528
rect 880 12848 17636 13128
rect 798 11768 17716 12848
rect 798 11488 17636 11768
rect 798 11088 17716 11488
rect 880 10808 17636 11088
rect 798 10408 17716 10808
rect 798 10128 17636 10408
rect 798 9728 17716 10128
rect 880 9448 17716 9728
rect 798 9048 17716 9448
rect 880 8768 17636 9048
rect 798 8368 17716 8768
rect 880 8088 17716 8368
rect 798 7688 17716 8088
rect 880 7408 17636 7688
rect 798 7008 17716 7408
rect 880 6728 17636 7008
rect 798 5648 17716 6728
rect 880 5368 17636 5648
rect 798 3608 17716 5368
rect 798 3328 17636 3608
rect 798 2928 17716 3328
rect 798 2648 17636 2928
rect 798 2143 17716 2648
<< metal4 >>
rect 2979 2128 3299 18000
rect 3639 2128 3959 18000
rect 7050 2128 7370 18000
rect 7710 2128 8030 18000
rect 11121 2128 11441 18000
rect 11781 2128 12101 18000
rect 15192 2128 15512 18000
rect 15852 2128 16172 18000
<< metal5 >>
rect 1056 16480 17436 16800
rect 1056 15820 17436 16140
rect 1056 12536 17436 12856
rect 1056 11876 17436 12196
rect 1056 8592 17436 8912
rect 1056 7932 17436 8252
rect 1056 4648 17436 4968
rect 1056 3988 17436 4308
<< labels >>
rlabel metal4 s 3639 2128 3959 18000 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 7710 2128 8030 18000 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 11781 2128 12101 18000 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 15852 2128 16172 18000 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 4648 17436 4968 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 8592 17436 8912 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 12536 17436 12856 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 16480 17436 16800 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 2979 2128 3299 18000 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 7050 2128 7370 18000 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 11121 2128 11441 18000 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 15192 2128 15512 18000 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 3988 17436 4308 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 7932 17436 8252 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 11876 17436 12196 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 15820 17436 16140 6 VPWR
port 2 nsew power bidirectional
rlabel metal3 s 17716 14288 18516 14408 6 a[0]
port 3 nsew signal input
rlabel metal2 s 5170 19860 5226 20660 6 a[10]
port 4 nsew signal input
rlabel metal3 s 0 15648 800 15768 6 a[11]
port 5 nsew signal input
rlabel metal2 s 10966 19860 11022 20660 6 a[12]
port 6 nsew signal input
rlabel metal2 s 9678 19860 9734 20660 6 a[13]
port 7 nsew signal input
rlabel metal2 s 12254 19860 12310 20660 6 a[14]
port 8 nsew signal input
rlabel metal2 s 8390 19860 8446 20660 6 a[15]
port 9 nsew signal input
rlabel metal3 s 0 12928 800 13048 6 a[16]
port 10 nsew signal input
rlabel metal3 s 0 13608 800 13728 6 a[17]
port 11 nsew signal input
rlabel metal3 s 0 10888 800 11008 6 a[18]
port 12 nsew signal input
rlabel metal3 s 0 9528 800 9648 6 a[19]
port 13 nsew signal input
rlabel metal3 s 17716 10888 18516 11008 6 a[1]
port 14 nsew signal input
rlabel metal3 s 0 8168 800 8288 6 a[20]
port 15 nsew signal input
rlabel metal2 s 8390 0 8446 800 6 a[21]
port 16 nsew signal input
rlabel metal2 s 5170 0 5226 800 6 a[22]
port 17 nsew signal input
rlabel metal2 s 9678 0 9734 800 6 a[23]
port 18 nsew signal input
rlabel metal2 s 12898 0 12954 800 6 a[24]
port 19 nsew signal input
rlabel metal3 s 17716 3408 18516 3528 6 a[25]
port 20 nsew signal input
rlabel metal3 s 17716 6808 18516 6928 6 a[26]
port 21 nsew signal input
rlabel metal3 s 17716 5448 18516 5568 6 a[27]
port 22 nsew signal input
rlabel metal2 s 10966 0 11022 800 6 a[28]
port 23 nsew signal input
rlabel metal2 s 7102 0 7158 800 6 a[29]
port 24 nsew signal input
rlabel metal3 s 17716 12928 18516 13048 6 a[2]
port 25 nsew signal input
rlabel metal3 s 0 5448 800 5568 6 a[30]
port 26 nsew signal input
rlabel metal3 s 0 7488 800 7608 6 a[31]
port 27 nsew signal input
rlabel metal3 s 17716 10208 18516 10328 6 a[3]
port 28 nsew signal input
rlabel metal3 s 17716 11568 18516 11688 6 a[4]
port 29 nsew signal input
rlabel metal3 s 17716 8848 18516 8968 6 a[5]
port 30 nsew signal input
rlabel metal3 s 17716 7488 18516 7608 6 a[6]
port 31 nsew signal input
rlabel metal2 s 10322 0 10378 800 6 a[7]
port 32 nsew signal input
rlabel metal3 s 0 8848 800 8968 6 a[8]
port 33 nsew signal input
rlabel metal2 s 9034 19860 9090 20660 6 a[9]
port 34 nsew signal input
rlabel metal3 s 0 17008 800 17128 6 clk
port 35 nsew signal input
rlabel metal3 s 17716 2728 18516 2848 6 rst
port 36 nsew signal input
rlabel metal3 s 0 6808 800 6928 6 x
port 37 nsew signal input
rlabel metal3 s 17716 14968 18516 15088 6 y
port 38 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 18516 20660
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 819092
string GDS_FILE /openlane/designs/spm/runs/run3/results/signoff/spm.magic.gds
string GDS_START 108486
<< end >>

