* NGSPICE file created from spm.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

.subckt spm VGND VPWR a[0] a[10] a[11] a[12] a[13] a[14] a[15] a[16] a[17] a[18] a[19]
+ a[1] a[20] a[21] a[22] a[23] a[24] a[25] a[26] a[27] a[28] a[29] a[2] a[30] a[31]
+ a[3] a[4] a[5] a[6] a[7] a[8] a[9] clk rst x y
X_294_ net47 dsa\[13\].last_carry_next net38 VGND VGND VPWR VPWR dsa\[13\].last_carry
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_15_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_12_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_277_ net50 dsa\[4\].y_out_next net41 VGND VGND VPWR VPWR dsa\[4\].y_out sky130_fd_sc_hd__dfrtp_1
X_200_ dsa\[19\].y_out _008_ _010_ VGND VGND VPWR VPWR dsa\[20\].last_carry_next sky130_fd_sc_hd__a21bo_1
X_131_ dsa\[5\].y_out _052_ VGND VGND VPWR VPWR dsa\[6\].y_out_next sky130_fd_sc_hd__xnor2_1
XFILLER_0_28_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_329_ net52 dsa\[30\].y_out_next net43 VGND VGND VPWR VPWR dsa\[30\].y_out sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_114_ _037_ _039_ VGND VGND VPWR VPWR _040_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_5_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_18_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_293_ net47 dsa\[12\].y_out_next net38 VGND VGND VPWR VPWR dsa\[12\].y_out sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_12_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_276_ net49 dsa\[4\].last_carry_next net40 VGND VGND VPWR VPWR dsa\[4\].last_carry
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_21_Right_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_130_ _050_ _051_ VGND VGND VPWR VPWR _052_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_72 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_259_ dsa\[15\].y_out _023_ VGND VGND VPWR VPWR dsa\[16\].y_out_next sky130_fd_sc_hd__xnor2_1
X_328_ net52 dsa\[30\].last_carry_next net43 VGND VGND VPWR VPWR dsa\[30\].last_carry
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_113_ _038_ net16 dsa\[8\].last_carry VGND VGND VPWR VPWR _039_ sky130_fd_sc_hd__nand3_1
XPHY_EDGE_ROW_8_Left_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_151 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_30 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_18_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_23_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_15_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_292_ net45 dsa\[12\].last_carry_next net36 VGND VGND VPWR VPWR dsa\[12\].last_carry
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_20_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_275_ net49 dsa\[3\].y_out_next net40 VGND VGND VPWR VPWR dsa\[3\].y_out sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_24_Left_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_258_ _021_ _022_ VGND VGND VPWR VPWR _023_ sky130_fd_sc_hd__nand2_1
X_327_ net52 dsa\[29\].y_out_next net43 VGND VGND VPWR VPWR dsa\[29\].y_out sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_189_ dsa\[0\].last_carry_next _095_ VGND VGND VPWR VPWR dsa\[0\].y_out_next sky130_fd_sc_hd__nor2_1
XFILLER_0_10_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_112_ _000_ VGND VGND VPWR VPWR _038_ sky130_fd_sc_hd__buf_2
XFILLER_0_24_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_11_Left_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_18_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_23_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_291_ net45 dsa\[11\].y_out_next net36 VGND VGND VPWR VPWR dsa\[11\].y_out sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_20_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_274_ net49 dsa\[3\].last_carry_next net40 VGND VGND VPWR VPWR dsa\[3\].last_carry
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_257_ _009_ net7 dsa\[16\].last_carry VGND VGND VPWR VPWR _022_ sky130_fd_sc_hd__nand3_1
X_326_ net51 dsa\[29\].last_carry_next net42 VGND VGND VPWR VPWR dsa\[29\].last_carry
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_188_ _009_ net25 dsa\[0\].last_carry VGND VGND VPWR VPWR _095_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_9_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_309_ net47 dsa\[20\].y_out_next net38 VGND VGND VPWR VPWR dsa\[20\].y_out sky130_fd_sc_hd__dfrtp_1
X_111_ _030_ net16 dsa\[8\].last_carry VGND VGND VPWR VPWR _037_ sky130_fd_sc_hd__a21o_1
XFILLER_0_15_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_6_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_290_ net45 dsa\[11\].last_carry_next net36 VGND VGND VPWR VPWR dsa\[11\].last_carry
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_3_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_273_ net46 dsa\[2\].y_out_next net37 VGND VGND VPWR VPWR dsa\[2\].y_out sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_256_ _001_ net7 dsa\[16\].last_carry VGND VGND VPWR VPWR _021_ sky130_fd_sc_hd__a21o_1
XFILLER_0_19_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_325_ net51 dsa\[28\].y_out_next net42 VGND VGND VPWR VPWR dsa\[28\].y_out sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_0_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_187_ _094_ VGND VGND VPWR VPWR dsa\[0\].last_carry_next sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_110_ dsa\[23\].y_out _036_ VGND VGND VPWR VPWR dsa\[24\].y_out_next sky130_fd_sc_hd__xnor2_1
XFILLER_0_27_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_308_ net47 dsa\[20\].last_carry_next net38 VGND VGND VPWR VPWR dsa\[20\].last_carry
+ sky130_fd_sc_hd__dfrtp_1
X_239_ _001_ net3 dsa\[20\].last_carry VGND VGND VPWR VPWR _008_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_10_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_6_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput35 net35 VGND VGND VPWR VPWR y sky130_fd_sc_hd__buf_2
XFILLER_0_7_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_28_Right_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_19_Right_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_272_ net45 dsa\[2\].last_carry_next net36 VGND VGND VPWR VPWR dsa\[2\].last_carry
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_255_ dsa\[17\].y_out _020_ VGND VGND VPWR VPWR dsa\[18\].y_out_next sky130_fd_sc_hd__xnor2_1
X_324_ net49 dsa\[28\].last_carry_next net40 VGND VGND VPWR VPWR dsa\[28\].last_carry
+ sky130_fd_sc_hd__dfrtp_1
X_186_ _000_ net25 dsa\[0\].last_carry VGND VGND VPWR VPWR _094_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_0_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_28_Left_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_307_ net47 dsa\[19\].y_out_next net38 VGND VGND VPWR VPWR dsa\[19\].y_out sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_238_ dsa\[1\].y_out _007_ VGND VGND VPWR VPWR dsa\[2\].y_out_next sky130_fd_sc_hd__xnor2_1
X_169_ dsa\[10\].y_out _081_ VGND VGND VPWR VPWR dsa\[11\].y_out_next sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_10_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_15_Left_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_3_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_24 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_0_Left_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_56 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_271_ net45 dsa\[1\].y_out_next net36 VGND VGND VPWR VPWR dsa\[1\].y_out sky130_fd_sc_hd__dfrtp_1
X_254_ _018_ _019_ VGND VGND VPWR VPWR _020_ sky130_fd_sc_hd__nand2_1
X_185_ dsa\[16\].y_out _093_ VGND VGND VPWR VPWR dsa\[17\].y_out_next sky130_fd_sc_hd__xnor2_1
X_323_ net51 dsa\[27\].y_out_next net42 VGND VGND VPWR VPWR dsa\[27\].y_out sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_306_ net51 dsa\[19\].last_carry_next net42 VGND VGND VPWR VPWR dsa\[19\].last_carry
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_3_Left_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_237_ _005_ _006_ VGND VGND VPWR VPWR _007_ sky130_fd_sc_hd__nand2_1
X_168_ _079_ _080_ VGND VGND VPWR VPWR _081_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_10_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_36 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_270_ net45 dsa\[1\].last_carry_next net36 VGND VGND VPWR VPWR dsa\[1\].last_carry
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_322_ net51 dsa\[27\].last_carry_next net42 VGND VGND VPWR VPWR dsa\[27\].last_carry
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_253_ _009_ net5 dsa\[18\].last_carry VGND VGND VPWR VPWR _019_ sky130_fd_sc_hd__nand3_1
X_184_ _091_ _092_ VGND VGND VPWR VPWR _093_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_0_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout50 net53 VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_18_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_305_ net51 dsa\[18\].y_out_next net42 VGND VGND VPWR VPWR dsa\[18\].y_out sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_236_ net22 _001_ dsa\[2\].last_carry VGND VGND VPWR VPWR _006_ sky130_fd_sc_hd__nand3_1
X_167_ _070_ net13 dsa\[11\].last_carry VGND VGND VPWR VPWR _080_ sky130_fd_sc_hd__nand3_1
XFILLER_0_15_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_219_ dsa\[26\].y_out _069_ _071_ VGND VGND VPWR VPWR dsa\[27\].last_carry_next sky130_fd_sc_hd__a21bo_1
XFILLER_0_27_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_24_Right_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_14_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout51 net53 VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__clkbuf_2
X_252_ _001_ net5 dsa\[18\].last_carry VGND VGND VPWR VPWR _018_ sky130_fd_sc_hd__a21o_1
X_183_ _070_ net6 dsa\[17\].last_carry VGND VGND VPWR VPWR _092_ sky130_fd_sc_hd__nand3_1
X_321_ net51 dsa\[26\].y_out_next net42 VGND VGND VPWR VPWR dsa\[26\].y_out sky130_fd_sc_hd__dfrtp_1
Xfanout40 net44 VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_304_ net48 dsa\[18\].last_carry_next net39 VGND VGND VPWR VPWR dsa\[18\].last_carry
+ sky130_fd_sc_hd__dfrtp_1
X_235_ net22 _000_ dsa\[2\].last_carry VGND VGND VPWR VPWR _005_ sky130_fd_sc_hd__a21o_1
XFILLER_0_24_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_166_ _062_ net13 dsa\[11\].last_carry VGND VGND VPWR VPWR _079_ sky130_fd_sc_hd__a21o_1
X_218_ dsa\[2\].y_out _066_ _067_ VGND VGND VPWR VPWR dsa\[3\].last_carry_next sky130_fd_sc_hd__a21bo_1
X_149_ _062_ net21 dsa\[3\].last_carry VGND VGND VPWR VPWR _066_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_17_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_19_Left_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout52 net53 VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__buf_1
X_182_ _062_ net6 dsa\[17\].last_carry VGND VGND VPWR VPWR _091_ sky130_fd_sc_hd__a21o_1
Xfanout41 net44 VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__buf_2
X_251_ dsa\[0\].y_out _017_ VGND VGND VPWR VPWR dsa\[1\].y_out_next sky130_fd_sc_hd__xnor2_1
X_320_ net50 dsa\[26\].last_carry_next net41 VGND VGND VPWR VPWR dsa\[26\].last_carry
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_303_ net51 dsa\[17\].y_out_next net42 VGND VGND VPWR VPWR dsa\[17\].y_out sky130_fd_sc_hd__dfrtp_1
X_165_ dsa\[28\].y_out _078_ VGND VGND VPWR VPWR dsa\[29\].y_out_next sky130_fd_sc_hd__xnor2_1
X_234_ dsa\[8\].y_out _004_ VGND VGND VPWR VPWR dsa\[9\].y_out_next sky130_fd_sc_hd__xnor2_1
XFILLER_0_1_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_7_Left_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_148_ dsa\[3\].y_out _065_ VGND VGND VPWR VPWR dsa\[4\].y_out_next sky130_fd_sc_hd__xnor2_1
X_217_ dsa\[3\].y_out _063_ _064_ VGND VGND VPWR VPWR dsa\[4\].last_carry_next sky130_fd_sc_hd__a21bo_1
XFILLER_0_12_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_17_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_20_Left_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout53 net33 VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__buf_2
X_181_ dsa\[21\].y_out _090_ VGND VGND VPWR VPWR dsa\[22\].y_out_next sky130_fd_sc_hd__xnor2_1
Xfanout42 net44 VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__clkbuf_4
X_250_ _015_ _016_ VGND VGND VPWR VPWR _017_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_302_ net51 dsa\[17\].last_carry_next net42 VGND VGND VPWR VPWR dsa\[17\].last_carry
+ sky130_fd_sc_hd__dfrtp_1
X_164_ _076_ _077_ VGND VGND VPWR VPWR _078_ sky130_fd_sc_hd__nand2_1
X_233_ _002_ _003_ VGND VGND VPWR VPWR _004_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_23_Left_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_61 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_147_ _063_ _064_ VGND VGND VPWR VPWR _065_ sky130_fd_sc_hd__nand2_1
X_216_ dsa\[25\].y_out _059_ _060_ VGND VGND VPWR VPWR dsa\[26\].last_carry_next sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_17_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_20_Right_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_180_ _088_ _089_ VGND VGND VPWR VPWR _090_ sky130_fd_sc_hd__nand2_1
Xfanout43 net44 VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_27_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_301_ net51 dsa\[16\].y_out_next net42 VGND VGND VPWR VPWR dsa\[16\].y_out sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_18 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_163_ _070_ net23 dsa\[29\].last_carry VGND VGND VPWR VPWR _077_ sky130_fd_sc_hd__nand3_1
X_232_ dsa\[9\].last_carry _001_ net15 VGND VGND VPWR VPWR _003_ sky130_fd_sc_hd__nand3_1
XFILLER_0_11_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_146_ _038_ net20 dsa\[4\].last_carry VGND VGND VPWR VPWR _064_ sky130_fd_sc_hd__nand3_1
X_215_ dsa\[4\].y_out _056_ _057_ VGND VGND VPWR VPWR dsa\[5\].last_carry_next sky130_fd_sc_hd__a21bo_1
XFILLER_0_12_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_72 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_129_ _038_ net18 dsa\[6\].last_carry VGND VGND VPWR VPWR _051_ sky130_fd_sc_hd__nand3_1
XFILLER_0_0_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout44 net34 VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__buf_2
XFILLER_0_3_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_300_ net48 dsa\[16\].last_carry_next net39 VGND VGND VPWR VPWR dsa\[16\].last_carry
+ sky130_fd_sc_hd__dfrtp_1
X_162_ _062_ net23 dsa\[29\].last_carry VGND VGND VPWR VPWR _076_ sky130_fd_sc_hd__a21o_1
X_231_ _001_ net15 dsa\[9\].last_carry VGND VGND VPWR VPWR _002_ sky130_fd_sc_hd__a21o_1
XFILLER_0_23_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput1 a[0] VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_214_ dsa\[27\].y_out _053_ _054_ VGND VGND VPWR VPWR dsa\[28\].last_carry_next sky130_fd_sc_hd__a21bo_1
X_145_ _062_ net20 dsa\[4\].last_carry VGND VGND VPWR VPWR _063_ sky130_fd_sc_hd__a21o_1
XFILLER_0_27_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_128_ _030_ net18 dsa\[6\].last_carry VGND VGND VPWR VPWR _050_ sky130_fd_sc_hd__a21o_1
XFILLER_0_7_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout45 net53 VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_25_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_161_ dsa\[30\].y_out _075_ VGND VGND VPWR VPWR dsa\[31\].y_out_next sky130_fd_sc_hd__xnor2_1
XFILLER_0_5_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_230_ _000_ VGND VGND VPWR VPWR _001_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_15_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput2 a[10] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_27_Left_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_213_ dsa\[5\].y_out _050_ _051_ VGND VGND VPWR VPWR dsa\[6\].last_carry_next sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_6_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_144_ _000_ VGND VGND VPWR VPWR _062_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_26_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_127_ dsa\[24\].y_out _049_ VGND VGND VPWR VPWR dsa\[25\].y_out_next sky130_fd_sc_hd__xnor2_1
XFILLER_0_21_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_14_Left_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout46 net53 VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_0_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_160_ _073_ _074_ VGND VGND VPWR VPWR _075_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_27_Right_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput3 a[11] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_18_Right_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_289_ net45 dsa\[10\].y_out_next net36 VGND VGND VPWR VPWR dsa\[10\].y_out sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_143_ dsa\[25\].y_out _061_ VGND VGND VPWR VPWR dsa\[26\].y_out_next sky130_fd_sc_hd__xnor2_1
XPHY_EDGE_ROW_2_Left_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_212_ dsa\[24\].y_out _047_ _048_ VGND VGND VPWR VPWR dsa\[25\].last_carry_next sky130_fd_sc_hd__a21bo_1
XFILLER_0_4_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_126_ _047_ _048_ VGND VGND VPWR VPWR _049_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_109_ _034_ _035_ VGND VGND VPWR VPWR _036_ sky130_fd_sc_hd__nand2_1
XFILLER_0_14_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout47 net53 VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__clkbuf_2
Xfanout36 net44 VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_26_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput4 a[12] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__buf_1
X_288_ net46 dsa\[10\].last_carry_next net37 VGND VGND VPWR VPWR dsa\[10\].last_carry
+ sky130_fd_sc_hd__dfrtp_1
X_142_ _059_ _060_ VGND VGND VPWR VPWR _061_ sky130_fd_sc_hd__nand2_1
X_211_ dsa\[6\].y_out _044_ _045_ VGND VGND VPWR VPWR dsa\[7\].last_carry_next sky130_fd_sc_hd__a21bo_1
X_125_ _038_ net29 dsa\[25\].last_carry VGND VGND VPWR VPWR _048_ sky130_fd_sc_hd__nand3_1
XFILLER_0_17_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_108_ _009_ net30 dsa\[24\].last_carry VGND VGND VPWR VPWR _035_ sky130_fd_sc_hd__nand3_1
XFILLER_0_8_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xfanout48 net53 VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__buf_1
Xfanout37 net44 VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_26_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput5 a[13] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_287_ net46 dsa\[9\].y_out_next net37 VGND VGND VPWR VPWR dsa\[10\].y_in sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_28_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_114 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_210_ dsa\[29\].y_out _041_ _042_ VGND VGND VPWR VPWR dsa\[30\].last_carry_next sky130_fd_sc_hd__a21bo_1
XFILLER_0_7_119 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_141_ _038_ net28 dsa\[26\].last_carry VGND VGND VPWR VPWR _060_ sky130_fd_sc_hd__nand3_1
XFILLER_0_11_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_124_ _030_ net29 dsa\[25\].last_carry VGND VGND VPWR VPWR _047_ sky130_fd_sc_hd__a21o_1
Xinput30 a[7] VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_13_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_107_ _030_ net30 dsa\[24\].last_carry VGND VGND VPWR VPWR _034_ sky130_fd_sc_hd__a21o_1
XFILLER_0_8_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_18_Left_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout38 net44 VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_14_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout49 net53 VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_26_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_286_ net45 dsa\[9\].last_carry_next net36 VGND VGND VPWR VPWR dsa\[9\].last_carry
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_79 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput6 a[14] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_23_Right_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_140_ _030_ net28 dsa\[26\].last_carry VGND VGND VPWR VPWR _059_ sky130_fd_sc_hd__a21o_1
X_269_ net45 dsa\[0\].y_out_next net36 VGND VGND VPWR VPWR dsa\[0\].y_out sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_6_Left_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_16_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_123_ dsa\[6\].y_out _046_ VGND VGND VPWR VPWR dsa\[7\].y_out_next sky130_fd_sc_hd__xnor2_1
XFILLER_0_3_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_7_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput20 a[27] VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__clkbuf_1
Xinput31 a[8] VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__buf_1
XFILLER_0_28_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_106_ dsa\[10\].y_in _033_ VGND VGND VPWR VPWR dsa\[10\].y_out_next sky130_fd_sc_hd__xnor2_1
XFILLER_0_28_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout39 net44 VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_25_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_285_ net46 dsa\[8\].y_out_next net37 VGND VGND VPWR VPWR dsa\[8\].y_out sky130_fd_sc_hd__dfrtp_1
Xinput7 a[15] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_22_Left_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_199_ dsa\[1\].y_out _005_ _006_ VGND VGND VPWR VPWR dsa\[2\].last_carry_next sky130_fd_sc_hd__a21bo_1
X_268_ net45 dsa\[0\].last_carry_next net36 VGND VGND VPWR VPWR dsa\[0\].last_carry
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_16_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_122_ _044_ _045_ VGND VGND VPWR VPWR _046_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_7_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput32 a[9] VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__buf_1
Xinput10 a[18] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__buf_1
Xinput21 a[28] VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_105_ _031_ _032_ VGND VGND VPWR VPWR _033_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_4_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_284_ net46 dsa\[8\].last_carry_next net37 VGND VGND VPWR VPWR dsa\[8\].last_carry
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput8 a[16] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__buf_1
XFILLER_0_14_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_267_ dsa\[11\].y_out _029_ VGND VGND VPWR VPWR dsa\[12\].y_out_next sky130_fd_sc_hd__xnor2_1
X_198_ dsa\[8\].y_out _002_ _003_ VGND VGND VPWR VPWR dsa\[9\].last_carry_next sky130_fd_sc_hd__a21bo_1
XTAP_TAPCELL_ROW_19_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_121_ _038_ net17 dsa\[7\].last_carry VGND VGND VPWR VPWR _045_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_11_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput33 clk VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__clkbuf_1
Xinput22 a[29] VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_7_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_319_ net50 dsa\[25\].y_out_next net41 VGND VGND VPWR VPWR dsa\[25\].y_out sky130_fd_sc_hd__dfrtp_1
Xinput11 a[19] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_28_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_104_ _009_ net14 dsa\[10\].last_carry VGND VGND VPWR VPWR _032_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_4_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_80 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput9 a[17] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__clkbuf_1
X_283_ net49 dsa\[7\].y_out_next net40 VGND VGND VPWR VPWR dsa\[7\].y_out sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_1_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_197_ dsa\[22\].y_out _101_ VGND VGND VPWR VPWR dsa\[23\].y_out_next sky130_fd_sc_hd__xnor2_1
X_266_ _027_ _028_ VGND VGND VPWR VPWR _029_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_120_ _030_ net17 dsa\[7\].last_carry VGND VGND VPWR VPWR _044_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_11_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput23 a[2] VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput12 a[1] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__clkbuf_1
Xinput34 rst VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__clkbuf_1
X_249_ _009_ net24 dsa\[1\].last_carry VGND VGND VPWR VPWR _016_ sky130_fd_sc_hd__nand3_1
X_318_ net49 dsa\[25\].last_carry_next net40 VGND VGND VPWR VPWR dsa\[25\].last_carry
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_91 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_103_ _030_ net14 dsa\[10\].last_carry VGND VGND VPWR VPWR _031_ sky130_fd_sc_hd__a21o_1
XFILLER_0_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_282_ net49 dsa\[7\].last_carry_next net40 VGND VGND VPWR VPWR dsa\[7\].last_carry
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_1_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_196_ _099_ _100_ VGND VGND VPWR VPWR _101_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_265_ _009_ net11 dsa\[12\].last_carry VGND VGND VPWR VPWR _028_ sky130_fd_sc_hd__nand3_1
XTAP_TAPCELL_ROW_25_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_26_Left_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_179_ _070_ net32 dsa\[22\].last_carry VGND VGND VPWR VPWR _089_ sky130_fd_sc_hd__nand3_1
XFILLER_0_17_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xinput24 a[30] VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__clkbuf_1
X_248_ _001_ net24 dsa\[1\].last_carry VGND VGND VPWR VPWR _015_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_10_Left_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput13 a[20] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__buf_1
X_317_ net49 dsa\[24\].y_out_next net40 VGND VGND VPWR VPWR dsa\[24\].y_out sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_22_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_102_ _000_ VGND VGND VPWR VPWR _030_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_20_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_13_Left_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_114 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_281_ net50 dsa\[6\].y_out_next net41 VGND VGND VPWR VPWR dsa\[6\].y_out sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_28_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_195_ _070_ net31 dsa\[23\].last_carry VGND VGND VPWR VPWR _100_ sky130_fd_sc_hd__nand3_1
X_264_ _001_ net11 dsa\[12\].last_carry VGND VGND VPWR VPWR _027_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_25_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_247_ dsa\[20\].y_out _014_ VGND VGND VPWR VPWR dsa\[21\].y_out_next sky130_fd_sc_hd__xnor2_1
XFILLER_0_17_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput14 a[21] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__buf_1
XPHY_EDGE_ROW_1_Left_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput25 a[31] VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__clkbuf_1
X_316_ net49 dsa\[24\].last_carry_next net40 VGND VGND VPWR VPWR dsa\[24\].last_carry
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_22_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_178_ _062_ net32 dsa\[22\].last_carry VGND VGND VPWR VPWR _088_ sky130_fd_sc_hd__a21o_1
XFILLER_0_3_128 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_126 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_280_ net50 dsa\[6\].last_carry_next net41 VGND VGND VPWR VPWR dsa\[6\].last_carry
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_13_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_28_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_263_ dsa\[13\].y_out _026_ VGND VGND VPWR VPWR dsa\[14\].y_out_next sky130_fd_sc_hd__xnor2_1
X_194_ _000_ net31 dsa\[23\].last_carry VGND VGND VPWR VPWR _099_ sky130_fd_sc_hd__a21o_1
XFILLER_0_10_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_25_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_246_ _012_ _013_ VGND VGND VPWR VPWR _014_ sky130_fd_sc_hd__nand2_1
X_177_ dsa\[18\].y_out _087_ VGND VGND VPWR VPWR dsa\[19\].y_out_next sky130_fd_sc_hd__xnor2_1
Xinput26 a[3] VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__buf_1
X_315_ net49 dsa\[23\].y_out_next net40 VGND VGND VPWR VPWR dsa\[23\].y_out sky130_fd_sc_hd__dfrtp_1
Xinput15 a[22] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__clkbuf_1
X_229_ x VGND VGND VPWR VPWR _000_ sky130_fd_sc_hd__buf_2
XFILLER_0_18_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_26_Right_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_28_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_331_ net52 dsa\[31\].y_out_next net43 VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__dfrtp_1
X_262_ _024_ _025_ VGND VGND VPWR VPWR _026_ sky130_fd_sc_hd__nand2_1
X_193_ dsa\[12\].y_out _098_ VGND VGND VPWR VPWR dsa\[13\].y_out_next sky130_fd_sc_hd__xnor2_1
XFILLER_0_6_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_71 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_111 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_245_ _009_ net2 dsa\[21\].last_carry VGND VGND VPWR VPWR _013_ sky130_fd_sc_hd__nand3_1
X_176_ _085_ _086_ VGND VGND VPWR VPWR _087_ sky130_fd_sc_hd__nand2_1
Xinput27 a[4] VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__buf_1
Xinput16 a[23] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__clkbuf_1
X_314_ net46 dsa\[23\].last_carry_next net37 VGND VGND VPWR VPWR dsa\[23\].last_carry
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_159_ _070_ net1 dsa\[31\].last_carry VGND VGND VPWR VPWR _074_ sky130_fd_sc_hd__nand3_1
X_228_ dsa\[22\].y_out _099_ _100_ VGND VGND VPWR VPWR dsa\[23\].last_carry_next sky130_fd_sc_hd__a21bo_1
XFILLER_0_20_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_17_Left_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_28_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_330_ net52 dsa\[31\].last_carry_next net43 VGND VGND VPWR VPWR dsa\[31\].last_carry
+ sky130_fd_sc_hd__dfrtp_1
X_261_ _009_ net9 dsa\[14\].last_carry VGND VGND VPWR VPWR _025_ sky130_fd_sc_hd__nand3_1
X_192_ _096_ _097_ VGND VGND VPWR VPWR _098_ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_131 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_106 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_244_ _001_ net2 dsa\[21\].last_carry VGND VGND VPWR VPWR _012_ sky130_fd_sc_hd__a21o_1
X_175_ _070_ net4 dsa\[19\].last_carry VGND VGND VPWR VPWR _086_ sky130_fd_sc_hd__nand3_1
X_313_ net48 dsa\[22\].y_out_next net39 VGND VGND VPWR VPWR dsa\[22\].y_out sky130_fd_sc_hd__dfrtp_1
Xinput17 a[24] VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput28 a[5] VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_5_Left_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_158_ _062_ net1 dsa\[31\].last_carry VGND VGND VPWR VPWR _073_ sky130_fd_sc_hd__a21o_1
XFILLER_0_18_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_227_ dsa\[12\].y_out _096_ _097_ VGND VGND VPWR VPWR dsa\[13\].last_carry_next sky130_fd_sc_hd__a21bo_1
XFILLER_0_20_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_28_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_260_ _001_ net9 dsa\[14\].last_carry VGND VGND VPWR VPWR _024_ sky130_fd_sc_hd__a21o_1
XFILLER_0_13_143 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_191_ _070_ net10 dsa\[13\].last_carry VGND VGND VPWR VPWR _097_ sky130_fd_sc_hd__nand3_1
XFILLER_0_6_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_243_ dsa\[19\].y_out _011_ VGND VGND VPWR VPWR dsa\[20\].y_out_next sky130_fd_sc_hd__xnor2_1
X_174_ _062_ net4 dsa\[19\].last_carry VGND VGND VPWR VPWR _085_ sky130_fd_sc_hd__a21o_1
X_312_ net48 dsa\[22\].last_carry_next net39 VGND VGND VPWR VPWR dsa\[22\].last_carry
+ sky130_fd_sc_hd__dfrtp_1
Xinput18 a[25] VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__clkbuf_1
Xinput29 a[6] VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_21_Left_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_226_ dsa\[16\].y_out _091_ _092_ VGND VGND VPWR VPWR dsa\[17\].last_carry_next sky130_fd_sc_hd__a21bo_1
XFILLER_0_18_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_157_ dsa\[26\].y_out _072_ VGND VGND VPWR VPWR dsa\[27\].y_out_next sky130_fd_sc_hd__xnor2_1
X_209_ dsa\[7\].y_out _037_ _039_ VGND VGND VPWR VPWR dsa\[8\].last_carry_next sky130_fd_sc_hd__a21bo_1
XFILLER_0_0_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_22_Right_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_190_ _000_ net10 dsa\[13\].last_carry VGND VGND VPWR VPWR _096_ sky130_fd_sc_hd__a21o_1
XFILLER_0_8_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_311_ net48 dsa\[21\].y_out_next net39 VGND VGND VPWR VPWR dsa\[21\].y_out sky130_fd_sc_hd__dfrtp_1
X_242_ _008_ _010_ VGND VGND VPWR VPWR _011_ sky130_fd_sc_hd__nand2_1
X_173_ dsa\[14\].y_out _084_ VGND VGND VPWR VPWR dsa\[15\].y_out_next sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_16_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput19 a[26] VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__clkbuf_1
X_225_ dsa\[21\].y_out _088_ _089_ VGND VGND VPWR VPWR dsa\[22\].last_carry_next sky130_fd_sc_hd__a21bo_1
XFILLER_0_18_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_156_ _069_ _071_ VGND VGND VPWR VPWR _072_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_139_ dsa\[4\].y_out _058_ VGND VGND VPWR VPWR dsa\[5\].y_out_next sky130_fd_sc_hd__xnor2_1
X_208_ dsa\[23\].y_out _034_ _035_ VGND VGND VPWR VPWR dsa\[24\].last_carry_next sky130_fd_sc_hd__a21bo_1
XFILLER_0_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_19_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_310_ net47 dsa\[21\].last_carry_next net38 VGND VGND VPWR VPWR dsa\[21\].last_carry
+ sky130_fd_sc_hd__dfrtp_1
X_241_ _009_ net3 dsa\[20\].last_carry VGND VGND VPWR VPWR _010_ sky130_fd_sc_hd__nand3_1
XFILLER_0_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_172_ _082_ _083_ VGND VGND VPWR VPWR _084_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_21_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_224_ dsa\[18\].y_out _085_ _086_ VGND VGND VPWR VPWR dsa\[19\].last_carry_next sky130_fd_sc_hd__a21bo_1
X_155_ _070_ net27 dsa\[27\].last_carry VGND VGND VPWR VPWR _071_ sky130_fd_sc_hd__nand3_1
XFILLER_0_18_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_9_Left_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_138_ _056_ _057_ VGND VGND VPWR VPWR _058_ sky130_fd_sc_hd__nand2_1
X_207_ dsa\[10\].y_in _031_ _032_ VGND VGND VPWR VPWR dsa\[10\].last_carry_next sky130_fd_sc_hd__a21bo_1
XFILLER_0_28_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_171_ _070_ net8 dsa\[15\].last_carry VGND VGND VPWR VPWR _083_ sky130_fd_sc_hd__nand3_1
X_240_ _000_ VGND VGND VPWR VPWR _009_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_223_ dsa\[14\].y_out _082_ _083_ VGND VGND VPWR VPWR dsa\[15\].last_carry_next sky130_fd_sc_hd__a21bo_1
XPHY_EDGE_ROW_25_Left_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_154_ _000_ VGND VGND VPWR VPWR _070_ sky130_fd_sc_hd__buf_2
X_137_ _038_ net19 dsa\[5\].last_carry VGND VGND VPWR VPWR _057_ sky130_fd_sc_hd__nand3_1
X_206_ dsa\[11\].y_out _027_ _028_ VGND VGND VPWR VPWR dsa\[12\].last_carry_next sky130_fd_sc_hd__a21bo_1
XFILLER_0_28_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_12_Left_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_27_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_170_ _062_ net8 dsa\[15\].last_carry VGND VGND VPWR VPWR _082_ sky130_fd_sc_hd__a21o_1
XFILLER_0_23_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_299_ net48 dsa\[15\].y_out_next net39 VGND VGND VPWR VPWR dsa\[15\].y_out sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_21_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_153_ _062_ net27 dsa\[27\].last_carry VGND VGND VPWR VPWR _069_ sky130_fd_sc_hd__a21o_1
X_222_ dsa\[10\].y_out _079_ _080_ VGND VGND VPWR VPWR dsa\[11\].last_carry_next sky130_fd_sc_hd__a21bo_1
XFILLER_0_20_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_205_ dsa\[13\].y_out _024_ _025_ VGND VGND VPWR VPWR dsa\[14\].last_carry_next sky130_fd_sc_hd__a21bo_1
X_136_ _030_ net19 dsa\[5\].last_carry VGND VGND VPWR VPWR _056_ sky130_fd_sc_hd__a21o_1
XFILLER_0_28_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_99 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_119_ dsa\[29\].y_out _043_ VGND VGND VPWR VPWR dsa\[30\].y_out_next sky130_fd_sc_hd__xnor2_1
XFILLER_0_15_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_112 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_27_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_298_ net47 dsa\[15\].last_carry_next net38 VGND VGND VPWR VPWR dsa\[15\].last_carry
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_221_ dsa\[28\].y_out _076_ _077_ VGND VGND VPWR VPWR dsa\[29\].last_carry_next sky130_fd_sc_hd__a21bo_1
X_152_ dsa\[2\].y_out _068_ VGND VGND VPWR VPWR dsa\[3\].y_out_next sky130_fd_sc_hd__xnor2_1
X_204_ dsa\[15\].y_out _021_ _022_ VGND VGND VPWR VPWR dsa\[16\].last_carry_next sky130_fd_sc_hd__a21bo_1
XFILLER_0_28_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_135_ dsa\[27\].y_out _055_ VGND VGND VPWR VPWR dsa\[28\].y_out_next sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_118_ _041_ _042_ VGND VGND VPWR VPWR _043_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_27_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_297_ net47 dsa\[14\].y_out_next net38 VGND VGND VPWR VPWR dsa\[14\].y_out sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_220_ dsa\[30\].y_out _073_ _074_ VGND VGND VPWR VPWR dsa\[31\].last_carry_next sky130_fd_sc_hd__a21bo_1
X_151_ _066_ _067_ VGND VGND VPWR VPWR _068_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_8_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_203_ dsa\[17\].y_out _018_ _019_ VGND VGND VPWR VPWR dsa\[18\].last_carry_next sky130_fd_sc_hd__a21bo_1
XFILLER_0_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_134_ _053_ _054_ VGND VGND VPWR VPWR _055_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_117_ _038_ net12 dsa\[30\].last_carry VGND VGND VPWR VPWR _042_ sky130_fd_sc_hd__nand3_1
XFILLER_0_21_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_16_Left_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_36 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_296_ net47 dsa\[14\].last_carry_next net38 VGND VGND VPWR VPWR dsa\[14\].last_carry
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_150_ _038_ net21 dsa\[3\].last_carry VGND VGND VPWR VPWR _067_ sky130_fd_sc_hd__nand3_1
XPHY_EDGE_ROW_25_Right_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_49 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_279_ net50 dsa\[5\].y_out_next net41 VGND VGND VPWR VPWR dsa\[5\].y_out sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_8_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_133_ _038_ net26 dsa\[28\].last_carry VGND VGND VPWR VPWR _054_ sky130_fd_sc_hd__nand3_1
XPHY_EDGE_ROW_4_Left_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_202_ dsa\[0\].y_out _015_ _016_ VGND VGND VPWR VPWR dsa\[1\].last_carry_next sky130_fd_sc_hd__a21bo_1
XFILLER_0_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_116_ _030_ net12 dsa\[30\].last_carry VGND VGND VPWR VPWR _041_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_5_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_48 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_295_ net47 dsa\[13\].y_out_next net38 VGND VGND VPWR VPWR dsa\[13\].y_out sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_278_ net50 dsa\[5\].last_carry_next net41 VGND VGND VPWR VPWR dsa\[5\].last_carry
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_201_ dsa\[20\].y_out _012_ _013_ VGND VGND VPWR VPWR dsa\[21\].last_carry_next sky130_fd_sc_hd__a21bo_1
XFILLER_0_20_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_132_ _030_ net26 dsa\[28\].last_carry VGND VGND VPWR VPWR _053_ sky130_fd_sc_hd__a21o_1
XFILLER_0_28_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_115_ dsa\[7\].y_out _040_ VGND VGND VPWR VPWR dsa\[8\].y_out_next sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_5_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
.ends

