magic
tech sky130A
magscale 1 2
timestamp 1742716265
<< nwell >>
rect 1066 2159 18254 19078
<< obsli1 >>
rect 1104 2159 18216 19057
<< obsm1 >>
rect 934 2128 18294 19088
<< metal2 >>
rect 1122 20742 1178 21542
rect 1674 20742 1730 21542
rect 2226 20742 2282 21542
rect 2778 20742 2834 21542
rect 3330 20742 3386 21542
rect 3882 20742 3938 21542
rect 4434 20742 4490 21542
rect 4986 20742 5042 21542
rect 5538 20742 5594 21542
rect 6090 20742 6146 21542
rect 6642 20742 6698 21542
rect 7194 20742 7250 21542
rect 7746 20742 7802 21542
rect 8298 20742 8354 21542
rect 8850 20742 8906 21542
rect 9402 20742 9458 21542
rect 9954 20742 10010 21542
rect 10506 20742 10562 21542
rect 11058 20742 11114 21542
rect 11610 20742 11666 21542
rect 12162 20742 12218 21542
rect 12714 20742 12770 21542
rect 13266 20742 13322 21542
rect 13818 20742 13874 21542
rect 14370 20742 14426 21542
rect 14922 20742 14978 21542
rect 15474 20742 15530 21542
rect 16026 20742 16082 21542
rect 16578 20742 16634 21542
rect 17130 20742 17186 21542
rect 17682 20742 17738 21542
rect 18234 20742 18290 21542
rect 14462 0 14518 800
<< obsm2 >>
rect 938 20686 1066 20890
rect 1234 20686 1618 20890
rect 1786 20686 2170 20890
rect 2338 20686 2722 20890
rect 2890 20686 3274 20890
rect 3442 20686 3826 20890
rect 3994 20686 4378 20890
rect 4546 20686 4930 20890
rect 5098 20686 5482 20890
rect 5650 20686 6034 20890
rect 6202 20686 6586 20890
rect 6754 20686 7138 20890
rect 7306 20686 7690 20890
rect 7858 20686 8242 20890
rect 8410 20686 8794 20890
rect 8962 20686 9346 20890
rect 9514 20686 9898 20890
rect 10066 20686 10450 20890
rect 10618 20686 11002 20890
rect 11170 20686 11554 20890
rect 11722 20686 12106 20890
rect 12274 20686 12658 20890
rect 12826 20686 13210 20890
rect 13378 20686 13762 20890
rect 13930 20686 14314 20890
rect 14482 20686 14866 20890
rect 15034 20686 15418 20890
rect 15586 20686 15970 20890
rect 16138 20686 16522 20890
rect 16690 20686 17074 20890
rect 17242 20686 17626 20890
rect 17794 20686 18178 20890
rect 938 856 18288 20686
rect 938 800 14406 856
rect 14574 800 18288 856
<< metal3 >>
rect 0 15784 800 15904
rect 18598 10616 19398 10736
rect 0 5176 800 5296
<< obsm3 >>
rect 800 15984 18598 19073
rect 880 15704 18598 15984
rect 800 10816 18598 15704
rect 800 10536 18518 10816
rect 800 5376 18598 10536
rect 880 5096 18598 5376
rect 800 2143 18598 5096
<< metal4 >>
rect 1904 2128 2304 19088
rect 2644 2128 3044 19088
rect 7904 2128 8304 19088
rect 8644 2128 9044 19088
rect 13904 2128 14304 19088
rect 14644 2128 15044 19088
<< obsm4 >>
rect 16619 5747 16685 18053
<< metal5 >>
rect 1056 15716 18264 16116
rect 1056 14976 18264 15376
rect 1056 9716 18264 10116
rect 1056 8976 18264 9376
rect 1056 3716 18264 4116
rect 1056 2976 18264 3376
<< labels >>
rlabel metal4 s 2644 2128 3044 19088 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 8644 2128 9044 19088 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 14644 2128 15044 19088 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 3716 18264 4116 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 9716 18264 10116 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 15716 18264 16116 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 1904 2128 2304 19088 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 7904 2128 8304 19088 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 13904 2128 14304 19088 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 2976 18264 3376 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 8976 18264 9376 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 14976 18264 15376 6 VPWR
port 2 nsew power bidirectional
rlabel metal2 s 1122 20742 1178 21542 6 a[0]
port 3 nsew signal input
rlabel metal2 s 6642 20742 6698 21542 6 a[10]
port 4 nsew signal input
rlabel metal2 s 7194 20742 7250 21542 6 a[11]
port 5 nsew signal input
rlabel metal2 s 7746 20742 7802 21542 6 a[12]
port 6 nsew signal input
rlabel metal2 s 8298 20742 8354 21542 6 a[13]
port 7 nsew signal input
rlabel metal2 s 8850 20742 8906 21542 6 a[14]
port 8 nsew signal input
rlabel metal2 s 9402 20742 9458 21542 6 a[15]
port 9 nsew signal input
rlabel metal2 s 9954 20742 10010 21542 6 a[16]
port 10 nsew signal input
rlabel metal2 s 10506 20742 10562 21542 6 a[17]
port 11 nsew signal input
rlabel metal2 s 11058 20742 11114 21542 6 a[18]
port 12 nsew signal input
rlabel metal2 s 11610 20742 11666 21542 6 a[19]
port 13 nsew signal input
rlabel metal2 s 1674 20742 1730 21542 6 a[1]
port 14 nsew signal input
rlabel metal2 s 12162 20742 12218 21542 6 a[20]
port 15 nsew signal input
rlabel metal2 s 12714 20742 12770 21542 6 a[21]
port 16 nsew signal input
rlabel metal2 s 13266 20742 13322 21542 6 a[22]
port 17 nsew signal input
rlabel metal2 s 13818 20742 13874 21542 6 a[23]
port 18 nsew signal input
rlabel metal2 s 14370 20742 14426 21542 6 a[24]
port 19 nsew signal input
rlabel metal2 s 14922 20742 14978 21542 6 a[25]
port 20 nsew signal input
rlabel metal2 s 15474 20742 15530 21542 6 a[26]
port 21 nsew signal input
rlabel metal2 s 16026 20742 16082 21542 6 a[27]
port 22 nsew signal input
rlabel metal2 s 16578 20742 16634 21542 6 a[28]
port 23 nsew signal input
rlabel metal2 s 17130 20742 17186 21542 6 a[29]
port 24 nsew signal input
rlabel metal2 s 2226 20742 2282 21542 6 a[2]
port 25 nsew signal input
rlabel metal2 s 17682 20742 17738 21542 6 a[30]
port 26 nsew signal input
rlabel metal2 s 18234 20742 18290 21542 6 a[31]
port 27 nsew signal input
rlabel metal2 s 2778 20742 2834 21542 6 a[3]
port 28 nsew signal input
rlabel metal2 s 3330 20742 3386 21542 6 a[4]
port 29 nsew signal input
rlabel metal2 s 3882 20742 3938 21542 6 a[5]
port 30 nsew signal input
rlabel metal2 s 4434 20742 4490 21542 6 a[6]
port 31 nsew signal input
rlabel metal2 s 4986 20742 5042 21542 6 a[7]
port 32 nsew signal input
rlabel metal2 s 5538 20742 5594 21542 6 a[8]
port 33 nsew signal input
rlabel metal2 s 6090 20742 6146 21542 6 a[9]
port 34 nsew signal input
rlabel metal3 s 18598 10616 19398 10736 6 clk
port 35 nsew signal input
rlabel metal2 s 14462 0 14518 800 6 rst
port 36 nsew signal input
rlabel metal3 s 0 15784 800 15904 6 x
port 37 nsew signal input
rlabel metal3 s 0 5176 800 5296 6 y
port 38 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 19398 21542
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 845838
string GDS_FILE /openlane/designs/spm/runs/openlane_test/results/signoff/spm.magic.gds
string GDS_START 144978
<< end >>

